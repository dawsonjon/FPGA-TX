//name : main_1
//input : input_socket:16
//input : input_rs232_rx:16
//input : input_switches:16
//input : input_buttons:16
//output : output_socket:16
//output : output_rs232_tx:16
//output : output_leds:16
//source_file : /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c

///+============================================================================+
///|                                                                            |
///|                     This file was generated by Chips                       |
///|                                                                            |
///|                                  Chips                                     |
///|                                                                            |
///|                      http://github.com/dawsonjon/Chips-2.0                 |
///|                                                                            |
///|                                                             Python powered |
///+============================================================================+
module main_1(input_socket,input_rs232_rx,input_switches,input_buttons,input_socket_stb,input_rs232_rx_stb,input_switches_stb,input_buttons_stb,output_socket_ack,output_rs232_tx_ack,output_leds_ack,clk,rst,output_socket,output_rs232_tx,output_leds,output_socket_stb,output_rs232_tx_stb,output_leds_stb,input_socket_ack,input_rs232_rx_ack,input_switches_ack,input_buttons_ack,exception);
  integer file_count;
  parameter  stop = 3'd0,
  instruction_fetch = 3'd1,
  operand_fetch = 3'd2,
  execute = 3'd3,
  load = 3'd4,
  wait_state = 3'd5,
  read = 3'd6,
  write = 3'd7;
  input [31:0] input_socket;
  input [31:0] input_rs232_rx;
  input [31:0] input_switches;
  input [31:0] input_buttons;
  input input_socket_stb;
  input input_rs232_rx_stb;
  input input_switches_stb;
  input input_buttons_stb;
  input output_socket_ack;
  input output_rs232_tx_ack;
  input output_leds_ack;
  input clk;
  input rst;
  output [31:0] output_socket;
  output [31:0] output_rs232_tx;
  output [31:0] output_leds;
  output output_socket_stb;
  output output_rs232_tx_stb;
  output output_leds_stb;
  output input_socket_ack;
  output input_rs232_rx_ack;
  output input_switches_ack;
  output input_buttons_ack;
  reg [31:0] timer;
  reg [63:0] timer_clock;
  reg [15:0] program_counter;
  reg [15:0] program_counter_1;
  reg [15:0] program_counter_2;
  reg [44:0] instruction;
  reg [4:0] opcode_2;
  reg [3:0] a;
  reg [3:0] b;
  reg [3:0] z;
  reg write_enable;
  reg [3:0] address_a_2;
  reg [3:0] address_b_2;
  reg [3:0] address_z_2;
  reg [3:0] address_z_3;
  reg [31:0] load_data;
  reg [31:0] write_output;
  reg [31:0] write_value;
  reg [31:0] read_input;
  reg [15:0] literal_2;
  reg [31:0] a_hi;
  reg [31:0] b_hi;
  reg [31:0] a_lo;
  reg [31:0] b_lo;
  reg [63:0] long_result;
  reg [31:0] result;
  reg [15:0] address;
  reg [31:0] data_out;
  reg [31:0] data_in;
  reg [31:0] carry;
  reg [31:0] s_output_socket_stb;
  reg [31:0] s_output_rs232_tx_stb;
  reg [31:0] s_output_leds_stb;
  reg [31:0] s_output_socket;
  reg [31:0] s_output_rs232_tx;
  reg [31:0] s_output_leds;
  reg [31:0] s_input_socket_ack;
  reg [31:0] s_input_rs232_rx_ack;
  reg [31:0] s_input_switches_ack;
  reg [31:0] s_input_buttons_ack;
  reg [7:0] state;
  output reg exception;
  reg [28:0] instructions [6636:0];
  reg [31:0] memory [4096:0];
  reg [31:0] registers [15:0];
  wire [31:0] operand_a;
  wire [31:0] operand_b;
  wire [31:0] register_a;
  wire [31:0] register_b;
  wire [15:0] literal;
  wire [4:0] opcode;
  wire [3:0] address_a;
  wire [3:0] address_b;
  wire [3:0] address_z;
  wire [15:0] load_address;
  wire [15:0] store_address;
  wire [31:0] store_data;
  wire  store_enable;

  //////////////////////////////////////////////////////////////////////////////
  // INSTRUCTION INITIALIZATION                                                 
  //                                                                            
  // Initialise the contents of the instruction memory                          
  //
  // Intruction Set
  // ==============
  // 0 {'literal': True, 'op': 'literal'}
  // 1 {'literal': True, 'op': 'addl'}
  // 2 {'literal': False, 'op': 'store'}
  // 3 {'literal': True, 'op': 'call'}
  // 4 {'literal': False, 'op': 'stop'}
  // 5 {'literal': False, 'op': 'load'}
  // 6 {'literal': False, 'op': 'read'}
  // 7 {'literal': False, 'op': 'unsigned_greater'}
  // 8 {'literal': True, 'op': 'jmp_if_false'}
  // 9 {'literal': False, 'op': 'unsigned_shift_right'}
  // 10 {'literal': False, 'op': 'and'}
  // 11 {'literal': False, 'op': 'add'}
  // 12 {'literal': True, 'op': 'goto'}
  // 13 {'literal': False, 'op': 'equal'}
  // 14 {'literal': True, 'op': 'jmp_if_true'}
  // 15 {'literal': False, 'op': 'not_equal'}
  // 16 {'literal': False, 'op': 'or'}
  // 17 {'literal': False, 'op': 'write'}
  // 18 {'literal': False, 'op': 'not'}
  // 19 {'literal': False, 'op': 'return'}
  // 20 {'literal': False, 'op': 'unsigned_greater_equal'}
  // 21 {'literal': False, 'op': 'subtract'}
  // 22 {'literal': False, 'op': 'shift_left'}
  // Intructions
  // ===========
  
  initial
  begin
    instructions[0] = {5'd0, 4'd3, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 183 {'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 183, 'op': 'literal'}
    instructions[1] = {5'd0, 4'd4, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 183 {'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 183, 'op': 'literal'}
    instructions[2] = {5'd1, 4'd3, 4'd3, 16'd96};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 183 {'a': 3, 'literal': 96, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 183, 'op': 'addl'}
    instructions[3] = {5'd0, 4'd8, 4'd0, 16'd13};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135 {'literal': 13, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135, 'op': 'literal'}
    instructions[4] = {5'd0, 4'd2, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135 {'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135, 'op': 'literal'}
    instructions[5] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135, 'op': 'store'}
    instructions[6] = {5'd0, 4'd8, 4'd0, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135 {'literal': 10, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135, 'op': 'literal'}
    instructions[7] = {5'd0, 4'd2, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135 {'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135, 'op': 'literal'}
    instructions[8] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135, 'op': 'store'}
    instructions[9] = {5'd0, 4'd8, 4'd0, 16'd13};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135 {'literal': 13, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135, 'op': 'literal'}
    instructions[10] = {5'd0, 4'd2, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135 {'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135, 'op': 'literal'}
    instructions[11] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135, 'op': 'store'}
    instructions[12] = {5'd0, 4'd8, 4'd0, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135 {'literal': 10, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135, 'op': 'literal'}
    instructions[13] = {5'd0, 4'd2, 4'd0, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135 {'literal': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135, 'op': 'literal'}
    instructions[14] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135, 'op': 'store'}
    instructions[15] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135, 'op': 'literal'}
    instructions[16] = {5'd0, 4'd2, 4'd0, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135 {'literal': 4, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135, 'op': 'literal'}
    instructions[17] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135, 'op': 'store'}
    instructions[18] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 18 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 18, 'op': 'literal'}
    instructions[19] = {5'd0, 4'd2, 4'd0, 16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 18 {'literal': 5, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 18, 'op': 'literal'}
    instructions[20] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 18 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 18, 'op': 'store'}
    instructions[21] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 5 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 5, 'op': 'literal'}
    instructions[22] = {5'd0, 4'd2, 4'd0, 16'd7};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 5 {'literal': 7, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 5, 'op': 'literal'}
    instructions[23] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 5 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 5, 'op': 'store'}
    instructions[24] = {5'd0, 4'd8, 4'd0, 16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 25 {'literal': 5, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 25, 'op': 'literal'}
    instructions[25] = {5'd0, 4'd2, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 25 {'literal': 8, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 25, 'op': 'literal'}
    instructions[26] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 25 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 25, 'op': 'store'}
    instructions[27] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 4 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 4, 'op': 'literal'}
    instructions[28] = {5'd0, 4'd2, 4'd0, 16'd9};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 4 {'literal': 9, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 4, 'op': 'literal'}
    instructions[29] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 4 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 4, 'op': 'store'}
    instructions[30] = {5'd0, 4'd8, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 26 {'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 26, 'op': 'literal'}
    instructions[31] = {5'd0, 4'd2, 4'd0, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 26 {'literal': 10, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 26, 'op': 'literal'}
    instructions[32] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 26 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 26, 'op': 'store'}
    instructions[33] = {5'd0, 4'd8, 4'd0, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 24 {'literal': 4, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 24, 'op': 'literal'}
    instructions[34] = {5'd0, 4'd2, 4'd0, 16'd11};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 24 {'literal': 11, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 24, 'op': 'literal'}
    instructions[35] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 24 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 24, 'op': 'store'}
    instructions[36] = {5'd0, 4'd8, 4'd0, 16'd87};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 87, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[37] = {5'd0, 4'd2, 4'd0, 16'd12};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 12, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[38] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'store'}
    instructions[39] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[40] = {5'd0, 4'd2, 4'd0, 16'd13};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 13, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[41] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'store'}
    instructions[42] = {5'd0, 4'd8, 4'd0, 16'd108};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 108, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[43] = {5'd0, 4'd2, 4'd0, 16'd14};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 14, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[44] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'store'}
    instructions[45] = {5'd0, 4'd8, 4'd0, 16'd99};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 99, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[46] = {5'd0, 4'd2, 4'd0, 16'd15};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 15, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[47] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'store'}
    instructions[48] = {5'd0, 4'd8, 4'd0, 16'd111};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 111, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[49] = {5'd0, 4'd2, 4'd0, 16'd16};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 16, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[50] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'store'}
    instructions[51] = {5'd0, 4'd8, 4'd0, 16'd109};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 109, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[52] = {5'd0, 4'd2, 4'd0, 16'd17};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 17, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[53] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'store'}
    instructions[54] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[55] = {5'd0, 4'd2, 4'd0, 16'd18};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 18, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[56] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'store'}
    instructions[57] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[58] = {5'd0, 4'd2, 4'd0, 16'd19};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 19, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[59] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'store'}
    instructions[60] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[61] = {5'd0, 4'd2, 4'd0, 16'd20};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 20, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[62] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'store'}
    instructions[63] = {5'd0, 4'd8, 4'd0, 16'd111};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 111, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[64] = {5'd0, 4'd2, 4'd0, 16'd21};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 21, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[65] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'store'}
    instructions[66] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[67] = {5'd0, 4'd2, 4'd0, 16'd22};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 22, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[68] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'store'}
    instructions[69] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[70] = {5'd0, 4'd2, 4'd0, 16'd23};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 23, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[71] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'store'}
    instructions[72] = {5'd0, 4'd8, 4'd0, 16'd104};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 104, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[73] = {5'd0, 4'd2, 4'd0, 16'd24};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 24, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[74] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'store'}
    instructions[75] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[76] = {5'd0, 4'd2, 4'd0, 16'd25};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 25, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[77] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'store'}
    instructions[78] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[79] = {5'd0, 4'd2, 4'd0, 16'd26};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 26, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[80] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'store'}
    instructions[81] = {5'd0, 4'd8, 4'd0, 16'd65};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 65, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[82] = {5'd0, 4'd2, 4'd0, 16'd27};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 27, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[83] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'store'}
    instructions[84] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[85] = {5'd0, 4'd2, 4'd0, 16'd28};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 28, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[86] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'store'}
    instructions[87] = {5'd0, 4'd8, 4'd0, 16'd108};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 108, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[88] = {5'd0, 4'd2, 4'd0, 16'd29};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 29, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[89] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'store'}
    instructions[90] = {5'd0, 4'd8, 4'd0, 16'd121};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 121, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[91] = {5'd0, 4'd2, 4'd0, 16'd30};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 30, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[92] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'store'}
    instructions[93] = {5'd0, 4'd8, 4'd0, 16'd115};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 115, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[94] = {5'd0, 4'd2, 4'd0, 16'd31};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 31, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[95] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'store'}
    instructions[96] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[97] = {5'd0, 4'd2, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 32, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[98] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'store'}
    instructions[99] = {5'd0, 4'd8, 4'd0, 16'd67};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 67, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[100] = {5'd0, 4'd2, 4'd0, 16'd33};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 33, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[101] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'store'}
    instructions[102] = {5'd0, 4'd8, 4'd0, 16'd104};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 104, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[103] = {5'd0, 4'd2, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 34, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[104] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'store'}
    instructions[105] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[106] = {5'd0, 4'd2, 4'd0, 16'd35};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 35, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[107] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'store'}
    instructions[108] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[109] = {5'd0, 4'd2, 4'd0, 16'd36};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 36, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[110] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'store'}
    instructions[111] = {5'd0, 4'd8, 4'd0, 16'd115};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 115, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[112] = {5'd0, 4'd2, 4'd0, 16'd37};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 37, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[113] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'store'}
    instructions[114] = {5'd0, 4'd8, 4'd0, 16'd45};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 45, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[115] = {5'd0, 4'd2, 4'd0, 16'd38};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 38, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[116] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'store'}
    instructions[117] = {5'd0, 4'd8, 4'd0, 16'd50};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 50, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[118] = {5'd0, 4'd2, 4'd0, 16'd39};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 39, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[119] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'store'}
    instructions[120] = {5'd0, 4'd8, 4'd0, 16'd46};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 46, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[121] = {5'd0, 4'd2, 4'd0, 16'd40};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 40, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[122] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'store'}
    instructions[123] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[124] = {5'd0, 4'd2, 4'd0, 16'd41};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 41, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[125] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'store'}
    instructions[126] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[127] = {5'd0, 4'd2, 4'd0, 16'd42};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 42, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[128] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'store'}
    instructions[129] = {5'd0, 4'd8, 4'd0, 16'd100};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 100, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[130] = {5'd0, 4'd2, 4'd0, 16'd43};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 43, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[131] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'store'}
    instructions[132] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[133] = {5'd0, 4'd2, 4'd0, 16'd44};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 44, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[134] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'store'}
    instructions[135] = {5'd0, 4'd8, 4'd0, 16'd109};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 109, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[136] = {5'd0, 4'd2, 4'd0, 16'd45};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 45, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[137] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'store'}
    instructions[138] = {5'd0, 4'd8, 4'd0, 16'd111};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 111, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[139] = {5'd0, 4'd2, 4'd0, 16'd46};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 46, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[140] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'store'}
    instructions[141] = {5'd0, 4'd8, 4'd0, 16'd33};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 33, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[142] = {5'd0, 4'd2, 4'd0, 16'd47};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 47, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[143] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'store'}
    instructions[144] = {5'd0, 4'd8, 4'd0, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 10, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[145] = {5'd0, 4'd2, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 48, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[146] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'store'}
    instructions[147] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[148] = {5'd0, 4'd2, 4'd0, 16'd49};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 49, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[149] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'store'}
    instructions[150] = {5'd0, 4'd8, 4'd0, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 22 {'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 22, 'op': 'literal'}
    instructions[151] = {5'd0, 4'd2, 4'd0, 16'd50};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 22 {'literal': 50, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 22, 'op': 'literal'}
    instructions[152] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 22 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 22, 'op': 'store'}
    instructions[153] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 14 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 14, 'op': 'literal'}
    instructions[154] = {5'd0, 4'd2, 4'd0, 16'd51};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 14 {'literal': 51, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 14, 'op': 'literal'}
    instructions[155] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 14 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 14, 'op': 'store'}
    instructions[156] = {5'd0, 4'd8, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 21 {'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 21, 'op': 'literal'}
    instructions[157] = {5'd0, 4'd2, 4'd0, 16'd52};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 21 {'literal': 52, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 21, 'op': 'literal'}
    instructions[158] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 21 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 21, 'op': 'store'}
    instructions[159] = {5'd0, 4'd8, 4'd0, 16'd67};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 67, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[160] = {5'd0, 4'd2, 4'd0, 16'd54};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 54, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[161] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'store'}
    instructions[162] = {5'd0, 4'd8, 4'd0, 16'd111};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 111, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[163] = {5'd0, 4'd2, 4'd0, 16'd55};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 55, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[164] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'store'}
    instructions[165] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[166] = {5'd0, 4'd2, 4'd0, 16'd56};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 56, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[167] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'store'}
    instructions[168] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[169] = {5'd0, 4'd2, 4'd0, 16'd57};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 57, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[170] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'store'}
    instructions[171] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[172] = {5'd0, 4'd2, 4'd0, 16'd58};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 58, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[173] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'store'}
    instructions[174] = {5'd0, 4'd8, 4'd0, 16'd99};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 99, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[175] = {5'd0, 4'd2, 4'd0, 16'd59};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 59, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[176] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'store'}
    instructions[177] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[178] = {5'd0, 4'd2, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 60, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[179] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'store'}
    instructions[180] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[181] = {5'd0, 4'd2, 4'd0, 16'd61};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 61, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[182] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'store'}
    instructions[183] = {5'd0, 4'd8, 4'd0, 16'd121};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 121, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[184] = {5'd0, 4'd2, 4'd0, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 62, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[185] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'store'}
    instructions[186] = {5'd0, 4'd8, 4'd0, 16'd111};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 111, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[187] = {5'd0, 4'd2, 4'd0, 16'd63};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 63, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[188] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'store'}
    instructions[189] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[190] = {5'd0, 4'd2, 4'd0, 16'd64};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 64, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[191] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'store'}
    instructions[192] = {5'd0, 4'd8, 4'd0, 16'd114};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 114, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[193] = {5'd0, 4'd2, 4'd0, 16'd65};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 65, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[194] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'store'}
    instructions[195] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[196] = {5'd0, 4'd2, 4'd0, 16'd66};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 66, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[197] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'store'}
    instructions[198] = {5'd0, 4'd8, 4'd0, 16'd119};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 119, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[199] = {5'd0, 4'd2, 4'd0, 16'd67};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 67, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[200] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'store'}
    instructions[201] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[202] = {5'd0, 4'd2, 4'd0, 16'd68};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 68, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[203] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'store'}
    instructions[204] = {5'd0, 4'd8, 4'd0, 16'd98};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 98, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[205] = {5'd0, 4'd2, 4'd0, 16'd69};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 69, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[206] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'store'}
    instructions[207] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[208] = {5'd0, 4'd2, 4'd0, 16'd70};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 70, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[209] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'store'}
    instructions[210] = {5'd0, 4'd8, 4'd0, 16'd98};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 98, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[211] = {5'd0, 4'd2, 4'd0, 16'd71};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 71, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[212] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'store'}
    instructions[213] = {5'd0, 4'd8, 4'd0, 16'd114};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 114, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[214] = {5'd0, 4'd2, 4'd0, 16'd72};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 72, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[215] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'store'}
    instructions[216] = {5'd0, 4'd8, 4'd0, 16'd111};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 111, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[217] = {5'd0, 4'd2, 4'd0, 16'd73};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 73, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[218] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'store'}
    instructions[219] = {5'd0, 4'd8, 4'd0, 16'd119};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 119, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[220] = {5'd0, 4'd2, 4'd0, 16'd74};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 74, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[221] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'store'}
    instructions[222] = {5'd0, 4'd8, 4'd0, 16'd115};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 115, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[223] = {5'd0, 4'd2, 4'd0, 16'd75};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 75, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[224] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'store'}
    instructions[225] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[226] = {5'd0, 4'd2, 4'd0, 16'd76};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 76, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[227] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'store'}
    instructions[228] = {5'd0, 4'd8, 4'd0, 16'd114};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 114, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[229] = {5'd0, 4'd2, 4'd0, 16'd77};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 77, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[230] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'store'}
    instructions[231] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[232] = {5'd0, 4'd2, 4'd0, 16'd78};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 78, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[233] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'store'}
    instructions[234] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[235] = {5'd0, 4'd2, 4'd0, 16'd79};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 79, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[236] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'store'}
    instructions[237] = {5'd0, 4'd8, 4'd0, 16'd111};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 111, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[238] = {5'd0, 4'd2, 4'd0, 16'd80};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 80, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[239] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'store'}
    instructions[240] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[241] = {5'd0, 4'd2, 4'd0, 16'd81};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 81, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[242] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'store'}
    instructions[243] = {5'd0, 4'd8, 4'd0, 16'd49};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 49, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[244] = {5'd0, 4'd2, 4'd0, 16'd82};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 82, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[245] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'store'}
    instructions[246] = {5'd0, 4'd8, 4'd0, 16'd57};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 57, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[247] = {5'd0, 4'd2, 4'd0, 16'd83};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 83, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[248] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'store'}
    instructions[249] = {5'd0, 4'd8, 4'd0, 16'd50};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 50, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[250] = {5'd0, 4'd2, 4'd0, 16'd84};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 84, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[251] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'store'}
    instructions[252] = {5'd0, 4'd8, 4'd0, 16'd46};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 46, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[253] = {5'd0, 4'd2, 4'd0, 16'd85};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 85, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[254] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'store'}
    instructions[255] = {5'd0, 4'd8, 4'd0, 16'd49};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 49, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[256] = {5'd0, 4'd2, 4'd0, 16'd86};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 86, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[257] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'store'}
    instructions[258] = {5'd0, 4'd8, 4'd0, 16'd54};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 54, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[259] = {5'd0, 4'd2, 4'd0, 16'd87};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 87, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[260] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'store'}
    instructions[261] = {5'd0, 4'd8, 4'd0, 16'd56};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 56, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[262] = {5'd0, 4'd2, 4'd0, 16'd88};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 88, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[263] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'store'}
    instructions[264] = {5'd0, 4'd8, 4'd0, 16'd46};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 46, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[265] = {5'd0, 4'd2, 4'd0, 16'd89};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 89, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[266] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'store'}
    instructions[267] = {5'd0, 4'd8, 4'd0, 16'd49};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 49, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[268] = {5'd0, 4'd2, 4'd0, 16'd90};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 90, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[269] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'store'}
    instructions[270] = {5'd0, 4'd8, 4'd0, 16'd46};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 46, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[271] = {5'd0, 4'd2, 4'd0, 16'd91};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 91, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[272] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'store'}
    instructions[273] = {5'd0, 4'd8, 4'd0, 16'd49};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 49, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[274] = {5'd0, 4'd2, 4'd0, 16'd92};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 92, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[275] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'store'}
    instructions[276] = {5'd0, 4'd8, 4'd0, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 10, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[277] = {5'd0, 4'd2, 4'd0, 16'd93};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 93, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[278] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'store'}
    instructions[279] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[280] = {5'd0, 4'd2, 4'd0, 16'd94};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 94, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[281] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'store'}
    instructions[282] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 19 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 19, 'op': 'literal'}
    instructions[283] = {5'd0, 4'd2, 4'd0, 16'd95};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 19 {'literal': 95, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 19, 'op': 'literal'}
    instructions[284] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 19 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 19, 'op': 'store'}
    instructions[285] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 183 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 183, 'op': 'addl'}
    instructions[286] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 183 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 183, 'op': 'addl'}
    instructions[287] = {5'd3, 4'd6, 4'd0, 16'd289};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 183 {'z': 6, 'label': 289, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 183, 'op': 'call'}
    instructions[288] = {5'd4, 4'd0, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 183 {'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 183, 'op': 'stop'}
    instructions[289] = {5'd1, 4'd3, 4'd3, 16'd2428};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 49 {'a': 3, 'literal': 2428, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 49, 'op': 'addl'}
    instructions[290] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 56 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 56, 'op': 'literal'}
    instructions[291] = {5'd1, 4'd2, 4'd4, 16'd1464};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 56 {'a': 4, 'literal': 1464, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 56, 'op': 'addl'}
    instructions[292] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 56 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 56, 'op': 'store'}
    instructions[293] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 57 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 57, 'op': 'literal'}
    instructions[294] = {5'd1, 4'd2, 4'd4, 16'd1465};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 57 {'a': 4, 'literal': 1465, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 57, 'op': 'addl'}
    instructions[295] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 57 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 57, 'op': 'store'}
    instructions[296] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 58 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 58, 'op': 'literal'}
    instructions[297] = {5'd1, 4'd2, 4'd4, 16'd1466};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 58 {'a': 4, 'literal': 1466, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 58, 'op': 'addl'}
    instructions[298] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 58 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 58, 'op': 'store'}
    instructions[299] = {5'd0, 4'd8, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 60, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[300] = {5'd1, 4'd2, 4'd4, 16'd1469};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1469, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[301] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[302] = {5'd0, 4'd8, 4'd0, 16'd104};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 104, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[303] = {5'd1, 4'd2, 4'd4, 16'd1470};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1470, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[304] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[305] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[306] = {5'd1, 4'd2, 4'd4, 16'd1471};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1471, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[307] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[308] = {5'd0, 4'd8, 4'd0, 16'd109};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 109, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[309] = {5'd1, 4'd2, 4'd4, 16'd1472};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1472, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[310] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[311] = {5'd0, 4'd8, 4'd0, 16'd108};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 108, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[312] = {5'd1, 4'd2, 4'd4, 16'd1473};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1473, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[313] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[314] = {5'd0, 4'd8, 4'd0, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 62, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[315] = {5'd1, 4'd2, 4'd4, 16'd1474};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1474, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[316] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[317] = {5'd0, 4'd8, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 60, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[318] = {5'd1, 4'd2, 4'd4, 16'd1475};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1475, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[319] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[320] = {5'd0, 4'd8, 4'd0, 16'd104};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 104, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[321] = {5'd1, 4'd2, 4'd4, 16'd1476};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1476, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[322] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[323] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[324] = {5'd1, 4'd2, 4'd4, 16'd1477};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1477, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[325] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[326] = {5'd0, 4'd8, 4'd0, 16'd97};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 97, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[327] = {5'd1, 4'd2, 4'd4, 16'd1478};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1478, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[328] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[329] = {5'd0, 4'd8, 4'd0, 16'd100};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 100, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[330] = {5'd1, 4'd2, 4'd4, 16'd1479};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1479, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[331] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[332] = {5'd0, 4'd8, 4'd0, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 62, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[333] = {5'd1, 4'd2, 4'd4, 16'd1480};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1480, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[334] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[335] = {5'd0, 4'd8, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 60, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[336] = {5'd1, 4'd2, 4'd4, 16'd1481};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1481, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[337] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[338] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[339] = {5'd1, 4'd2, 4'd4, 16'd1482};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1482, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[340] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[341] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[342] = {5'd1, 4'd2, 4'd4, 16'd1483};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1483, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[343] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[344] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[345] = {5'd1, 4'd2, 4'd4, 16'd1484};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1484, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[346] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[347] = {5'd0, 4'd8, 4'd0, 16'd108};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 108, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[348] = {5'd1, 4'd2, 4'd4, 16'd1485};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1485, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[349] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[350] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[351] = {5'd1, 4'd2, 4'd4, 16'd1486};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1486, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[352] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[353] = {5'd0, 4'd8, 4'd0, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 62, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[354] = {5'd1, 4'd2, 4'd4, 16'd1487};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1487, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[355] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[356] = {5'd0, 4'd8, 4'd0, 16'd67};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 67, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[357] = {5'd1, 4'd2, 4'd4, 16'd1488};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1488, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[358] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[359] = {5'd0, 4'd8, 4'd0, 16'd104};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 104, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[360] = {5'd1, 4'd2, 4'd4, 16'd1489};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1489, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[361] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[362] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[363] = {5'd1, 4'd2, 4'd4, 16'd1490};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1490, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[364] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[365] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[366] = {5'd1, 4'd2, 4'd4, 16'd1491};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1491, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[367] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[368] = {5'd0, 4'd8, 4'd0, 16'd115};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 115, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[369] = {5'd1, 4'd2, 4'd4, 16'd1492};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1492, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[370] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[371] = {5'd0, 4'd8, 4'd0, 16'd45};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 45, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[372] = {5'd1, 4'd2, 4'd4, 16'd1493};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1493, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[373] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[374] = {5'd0, 4'd8, 4'd0, 16'd50};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 50, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[375] = {5'd1, 4'd2, 4'd4, 16'd1494};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1494, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[376] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[377] = {5'd0, 4'd8, 4'd0, 16'd46};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 46, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[378] = {5'd1, 4'd2, 4'd4, 16'd1495};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1495, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[379] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[380] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[381] = {5'd1, 4'd2, 4'd4, 16'd1496};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1496, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[382] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[383] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[384] = {5'd1, 4'd2, 4'd4, 16'd1497};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1497, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[385] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[386] = {5'd0, 4'd8, 4'd0, 16'd65};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 65, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[387] = {5'd1, 4'd2, 4'd4, 16'd1498};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1498, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[388] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[389] = {5'd0, 4'd8, 4'd0, 16'd84};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 84, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[390] = {5'd1, 4'd2, 4'd4, 16'd1499};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1499, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[391] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[392] = {5'd0, 4'd8, 4'd0, 16'd76};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 76, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[393] = {5'd1, 4'd2, 4'd4, 16'd1500};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1500, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[394] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[395] = {5'd0, 4'd8, 4'd0, 16'd89};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 89, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[396] = {5'd1, 4'd2, 4'd4, 16'd1501};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1501, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[397] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[398] = {5'd0, 4'd8, 4'd0, 16'd83};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 83, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[399] = {5'd1, 4'd2, 4'd4, 16'd1502};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1502, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[400] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[401] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[402] = {5'd1, 4'd2, 4'd4, 16'd1503};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1503, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[403] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[404] = {5'd0, 4'd8, 4'd0, 16'd68};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 68, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[405] = {5'd1, 4'd2, 4'd4, 16'd1504};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1504, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[406] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[407] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[408] = {5'd1, 4'd2, 4'd4, 16'd1505};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1505, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[409] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[410] = {5'd0, 4'd8, 4'd0, 16'd109};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 109, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[411] = {5'd1, 4'd2, 4'd4, 16'd1506};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1506, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[412] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[413] = {5'd0, 4'd8, 4'd0, 16'd111};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 111, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[414] = {5'd1, 4'd2, 4'd4, 16'd1507};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1507, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[415] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[416] = {5'd0, 4'd8, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 60, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[417] = {5'd1, 4'd2, 4'd4, 16'd1508};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1508, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[418] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[419] = {5'd0, 4'd8, 4'd0, 16'd47};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 47, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[420] = {5'd1, 4'd2, 4'd4, 16'd1509};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1509, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[421] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[422] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[423] = {5'd1, 4'd2, 4'd4, 16'd1510};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1510, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[424] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[425] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[426] = {5'd1, 4'd2, 4'd4, 16'd1511};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1511, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[427] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[428] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[429] = {5'd1, 4'd2, 4'd4, 16'd1512};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1512, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[430] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[431] = {5'd0, 4'd8, 4'd0, 16'd108};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 108, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[432] = {5'd1, 4'd2, 4'd4, 16'd1513};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1513, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[433] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[434] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[435] = {5'd1, 4'd2, 4'd4, 16'd1514};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1514, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[436] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[437] = {5'd0, 4'd8, 4'd0, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 62, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[438] = {5'd1, 4'd2, 4'd4, 16'd1515};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1515, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[439] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[440] = {5'd0, 4'd8, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 60, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[441] = {5'd1, 4'd2, 4'd4, 16'd1516};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1516, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[442] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[443] = {5'd0, 4'd8, 4'd0, 16'd47};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 47, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[444] = {5'd1, 4'd2, 4'd4, 16'd1517};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1517, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[445] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[446] = {5'd0, 4'd8, 4'd0, 16'd104};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 104, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[447] = {5'd1, 4'd2, 4'd4, 16'd1518};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1518, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[448] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[449] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[450] = {5'd1, 4'd2, 4'd4, 16'd1519};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1519, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[451] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[452] = {5'd0, 4'd8, 4'd0, 16'd97};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 97, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[453] = {5'd1, 4'd2, 4'd4, 16'd1520};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1520, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[454] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[455] = {5'd0, 4'd8, 4'd0, 16'd100};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 100, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[456] = {5'd1, 4'd2, 4'd4, 16'd1521};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1521, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[457] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[458] = {5'd0, 4'd8, 4'd0, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 62, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[459] = {5'd1, 4'd2, 4'd4, 16'd1522};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1522, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[460] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[461] = {5'd0, 4'd8, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 60, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[462] = {5'd1, 4'd2, 4'd4, 16'd1523};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1523, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[463] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[464] = {5'd0, 4'd8, 4'd0, 16'd98};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 98, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[465] = {5'd1, 4'd2, 4'd4, 16'd1524};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1524, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[466] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[467] = {5'd0, 4'd8, 4'd0, 16'd111};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 111, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[468] = {5'd1, 4'd2, 4'd4, 16'd1525};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1525, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[469] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[470] = {5'd0, 4'd8, 4'd0, 16'd100};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 100, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[471] = {5'd1, 4'd2, 4'd4, 16'd1526};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1526, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[472] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[473] = {5'd0, 4'd8, 4'd0, 16'd121};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 121, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[474] = {5'd1, 4'd2, 4'd4, 16'd1527};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1527, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[475] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[476] = {5'd0, 4'd8, 4'd0, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 62, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[477] = {5'd1, 4'd2, 4'd4, 16'd1528};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1528, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[478] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[479] = {5'd0, 4'd8, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 60, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[480] = {5'd1, 4'd2, 4'd4, 16'd1529};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1529, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[481] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[482] = {5'd0, 4'd8, 4'd0, 16'd104};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 104, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[483] = {5'd1, 4'd2, 4'd4, 16'd1530};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1530, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[484] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[485] = {5'd0, 4'd8, 4'd0, 16'd49};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 49, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[486] = {5'd1, 4'd2, 4'd4, 16'd1531};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1531, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[487] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[488] = {5'd0, 4'd8, 4'd0, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 62, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[489] = {5'd1, 4'd2, 4'd4, 16'd1532};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1532, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[490] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[491] = {5'd0, 4'd8, 4'd0, 16'd67};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 67, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[492] = {5'd1, 4'd2, 4'd4, 16'd1533};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1533, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[493] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[494] = {5'd0, 4'd8, 4'd0, 16'd104};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 104, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[495] = {5'd1, 4'd2, 4'd4, 16'd1534};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1534, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[496] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[497] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[498] = {5'd1, 4'd2, 4'd4, 16'd1535};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1535, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[499] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[500] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[501] = {5'd1, 4'd2, 4'd4, 16'd1536};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1536, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[502] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[503] = {5'd0, 4'd8, 4'd0, 16'd115};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 115, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[504] = {5'd1, 4'd2, 4'd4, 16'd1537};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1537, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[505] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[506] = {5'd0, 4'd8, 4'd0, 16'd45};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 45, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[507] = {5'd1, 4'd2, 4'd4, 16'd1538};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1538, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[508] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[509] = {5'd0, 4'd8, 4'd0, 16'd50};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 50, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[510] = {5'd1, 4'd2, 4'd4, 16'd1539};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1539, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[511] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[512] = {5'd0, 4'd8, 4'd0, 16'd46};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 46, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[513] = {5'd1, 4'd2, 4'd4, 16'd1540};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1540, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[514] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[515] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[516] = {5'd1, 4'd2, 4'd4, 16'd1541};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1541, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[517] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[518] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[519] = {5'd1, 4'd2, 4'd4, 16'd1542};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1542, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[520] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[521] = {5'd0, 4'd8, 4'd0, 16'd65};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 65, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[522] = {5'd1, 4'd2, 4'd4, 16'd1543};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1543, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[523] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[524] = {5'd0, 4'd8, 4'd0, 16'd84};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 84, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[525] = {5'd1, 4'd2, 4'd4, 16'd1544};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1544, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[526] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[527] = {5'd0, 4'd8, 4'd0, 16'd76};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 76, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[528] = {5'd1, 4'd2, 4'd4, 16'd1545};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1545, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[529] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[530] = {5'd0, 4'd8, 4'd0, 16'd89};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 89, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[531] = {5'd1, 4'd2, 4'd4, 16'd1546};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1546, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[532] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[533] = {5'd0, 4'd8, 4'd0, 16'd83};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 83, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[534] = {5'd1, 4'd2, 4'd4, 16'd1547};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1547, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[535] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[536] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[537] = {5'd1, 4'd2, 4'd4, 16'd1548};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1548, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[538] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[539] = {5'd0, 4'd8, 4'd0, 16'd68};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 68, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[540] = {5'd1, 4'd2, 4'd4, 16'd1549};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1549, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[541] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[542] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[543] = {5'd1, 4'd2, 4'd4, 16'd1550};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1550, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[544] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[545] = {5'd0, 4'd8, 4'd0, 16'd109};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 109, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[546] = {5'd1, 4'd2, 4'd4, 16'd1551};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1551, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[547] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[548] = {5'd0, 4'd8, 4'd0, 16'd111};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 111, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[549] = {5'd1, 4'd2, 4'd4, 16'd1552};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1552, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[550] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[551] = {5'd0, 4'd8, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 60, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[552] = {5'd1, 4'd2, 4'd4, 16'd1553};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1553, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[553] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[554] = {5'd0, 4'd8, 4'd0, 16'd47};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 47, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[555] = {5'd1, 4'd2, 4'd4, 16'd1554};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1554, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[556] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[557] = {5'd0, 4'd8, 4'd0, 16'd104};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 104, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[558] = {5'd1, 4'd2, 4'd4, 16'd1555};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1555, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[559] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[560] = {5'd0, 4'd8, 4'd0, 16'd49};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 49, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[561] = {5'd1, 4'd2, 4'd4, 16'd1556};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1556, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[562] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[563] = {5'd0, 4'd8, 4'd0, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 62, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[564] = {5'd1, 4'd2, 4'd4, 16'd1557};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1557, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[565] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[566] = {5'd0, 4'd8, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 60, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[567] = {5'd1, 4'd2, 4'd4, 16'd1558};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1558, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[568] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[569] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[570] = {5'd1, 4'd2, 4'd4, 16'd1559};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1559, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[571] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[572] = {5'd0, 4'd8, 4'd0, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 62, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[573] = {5'd1, 4'd2, 4'd4, 16'd1560};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1560, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[574] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[575] = {5'd0, 4'd8, 4'd0, 16'd87};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 87, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[576] = {5'd1, 4'd2, 4'd4, 16'd1561};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1561, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[577] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[578] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[579] = {5'd1, 4'd2, 4'd4, 16'd1562};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1562, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[580] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[581] = {5'd0, 4'd8, 4'd0, 16'd108};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 108, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[582] = {5'd1, 4'd2, 4'd4, 16'd1563};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1563, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[583] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[584] = {5'd0, 4'd8, 4'd0, 16'd99};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 99, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[585] = {5'd1, 4'd2, 4'd4, 16'd1564};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1564, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[586] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[587] = {5'd0, 4'd8, 4'd0, 16'd111};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 111, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[588] = {5'd1, 4'd2, 4'd4, 16'd1565};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1565, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[589] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[590] = {5'd0, 4'd8, 4'd0, 16'd109};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 109, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[591] = {5'd1, 4'd2, 4'd4, 16'd1566};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1566, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[592] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[593] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[594] = {5'd1, 4'd2, 4'd4, 16'd1567};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1567, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[595] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[596] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[597] = {5'd1, 4'd2, 4'd4, 16'd1568};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1568, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[598] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[599] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[600] = {5'd1, 4'd2, 4'd4, 16'd1569};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1569, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[601] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[602] = {5'd0, 4'd8, 4'd0, 16'd111};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 111, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[603] = {5'd1, 4'd2, 4'd4, 16'd1570};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1570, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[604] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[605] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[606] = {5'd1, 4'd2, 4'd4, 16'd1571};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1571, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[607] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[608] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[609] = {5'd1, 4'd2, 4'd4, 16'd1572};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1572, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[610] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[611] = {5'd0, 4'd8, 4'd0, 16'd104};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 104, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[612] = {5'd1, 4'd2, 4'd4, 16'd1573};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1573, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[613] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[614] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[615] = {5'd1, 4'd2, 4'd4, 16'd1574};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1574, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[616] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[617] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[618] = {5'd1, 4'd2, 4'd4, 16'd1575};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1575, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[619] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[620] = {5'd0, 4'd8, 4'd0, 16'd67};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 67, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[621] = {5'd1, 4'd2, 4'd4, 16'd1576};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1576, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[622] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[623] = {5'd0, 4'd8, 4'd0, 16'd104};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 104, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[624] = {5'd1, 4'd2, 4'd4, 16'd1577};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1577, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[625] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[626] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[627] = {5'd1, 4'd2, 4'd4, 16'd1578};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1578, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[628] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[629] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[630] = {5'd1, 4'd2, 4'd4, 16'd1579};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1579, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[631] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[632] = {5'd0, 4'd8, 4'd0, 16'd115};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 115, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[633] = {5'd1, 4'd2, 4'd4, 16'd1580};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1580, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[634] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[635] = {5'd0, 4'd8, 4'd0, 16'd45};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 45, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[636] = {5'd1, 4'd2, 4'd4, 16'd1581};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1581, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[637] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[638] = {5'd0, 4'd8, 4'd0, 16'd50};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 50, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[639] = {5'd1, 4'd2, 4'd4, 16'd1582};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1582, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[640] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[641] = {5'd0, 4'd8, 4'd0, 16'd46};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 46, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[642] = {5'd1, 4'd2, 4'd4, 16'd1583};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1583, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[643] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[644] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[645] = {5'd1, 4'd2, 4'd4, 16'd1584};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1584, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[646] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[647] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[648] = {5'd1, 4'd2, 4'd4, 16'd1585};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1585, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[649] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[650] = {5'd0, 4'd8, 4'd0, 16'd65};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 65, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[651] = {5'd1, 4'd2, 4'd4, 16'd1586};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1586, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[652] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[653] = {5'd0, 4'd8, 4'd0, 16'd84};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 84, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[654] = {5'd1, 4'd2, 4'd4, 16'd1587};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1587, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[655] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[656] = {5'd0, 4'd8, 4'd0, 16'd76};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 76, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[657] = {5'd1, 4'd2, 4'd4, 16'd1588};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1588, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[658] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[659] = {5'd0, 4'd8, 4'd0, 16'd89};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 89, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[660] = {5'd1, 4'd2, 4'd4, 16'd1589};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1589, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[661] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[662] = {5'd0, 4'd8, 4'd0, 16'd83};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 83, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[663] = {5'd1, 4'd2, 4'd4, 16'd1590};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1590, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[664] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[665] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[666] = {5'd1, 4'd2, 4'd4, 16'd1591};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1591, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[667] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[668] = {5'd0, 4'd8, 4'd0, 16'd68};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 68, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[669] = {5'd1, 4'd2, 4'd4, 16'd1592};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1592, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[670] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[671] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[672] = {5'd1, 4'd2, 4'd4, 16'd1593};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1593, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[673] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[674] = {5'd0, 4'd8, 4'd0, 16'd109};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 109, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[675] = {5'd1, 4'd2, 4'd4, 16'd1594};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1594, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[676] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[677] = {5'd0, 4'd8, 4'd0, 16'd111};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 111, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[678] = {5'd1, 4'd2, 4'd4, 16'd1595};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1595, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[679] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[680] = {5'd0, 4'd8, 4'd0, 16'd33};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 33, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[681] = {5'd1, 4'd2, 4'd4, 16'd1596};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1596, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[682] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[683] = {5'd0, 4'd8, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 60, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[684] = {5'd1, 4'd2, 4'd4, 16'd1597};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1597, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[685] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[686] = {5'd0, 4'd8, 4'd0, 16'd47};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 47, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[687] = {5'd1, 4'd2, 4'd4, 16'd1598};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1598, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[688] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[689] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[690] = {5'd1, 4'd2, 4'd4, 16'd1599};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1599, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[691] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[692] = {5'd0, 4'd8, 4'd0, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 62, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[693] = {5'd1, 4'd2, 4'd4, 16'd1600};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1600, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[694] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[695] = {5'd0, 4'd8, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 60, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[696] = {5'd1, 4'd2, 4'd4, 16'd1601};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1601, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[697] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[698] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[699] = {5'd1, 4'd2, 4'd4, 16'd1602};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1602, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[700] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[701] = {5'd0, 4'd8, 4'd0, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 62, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[702] = {5'd1, 4'd2, 4'd4, 16'd1603};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1603, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[703] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[704] = {5'd0, 4'd8, 4'd0, 16'd83};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 83, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[705] = {5'd1, 4'd2, 4'd4, 16'd1604};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1604, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[706] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[707] = {5'd0, 4'd8, 4'd0, 16'd119};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 119, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[708] = {5'd1, 4'd2, 4'd4, 16'd1605};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1605, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[709] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[710] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[711] = {5'd1, 4'd2, 4'd4, 16'd1606};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1606, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[712] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[713] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[714] = {5'd1, 4'd2, 4'd4, 16'd1607};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1607, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[715] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[716] = {5'd0, 4'd8, 4'd0, 16'd99};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 99, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[717] = {5'd1, 4'd2, 4'd4, 16'd1608};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1608, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[718] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[719] = {5'd0, 4'd8, 4'd0, 16'd104};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 104, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[720] = {5'd1, 4'd2, 4'd4, 16'd1609};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1609, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[721] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[722] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[723] = {5'd1, 4'd2, 4'd4, 16'd1610};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1610, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[724] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[725] = {5'd0, 4'd8, 4'd0, 16'd83};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 83, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[726] = {5'd1, 4'd2, 4'd4, 16'd1611};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1611, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[727] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[728] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[729] = {5'd1, 4'd2, 4'd4, 16'd1612};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1612, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[730] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[731] = {5'd0, 4'd8, 4'd0, 16'd97};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 97, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[732] = {5'd1, 4'd2, 4'd4, 16'd1613};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1613, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[733] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[734] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[735] = {5'd1, 4'd2, 4'd4, 16'd1614};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1614, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[736] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[737] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[738] = {5'd1, 4'd2, 4'd4, 16'd1615};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1615, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[739] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[740] = {5'd0, 4'd8, 4'd0, 16'd115};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 115, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[741] = {5'd1, 4'd2, 4'd4, 16'd1616};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1616, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[742] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[743] = {5'd0, 4'd8, 4'd0, 16'd58};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 58, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[744] = {5'd1, 4'd2, 4'd4, 16'd1617};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1617, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[745] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[746] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[747] = {5'd1, 4'd2, 4'd4, 16'd1618};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1618, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[748] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[749] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[750] = {5'd1, 4'd2, 4'd4, 16'd1619};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1619, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[751] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[752] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[753] = {5'd1, 4'd2, 4'd4, 16'd1620};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1620, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[754] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[755] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[756] = {5'd1, 4'd2, 4'd4, 16'd1621};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1621, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[757] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[758] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[759] = {5'd1, 4'd2, 4'd4, 16'd1622};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1622, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[760] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[761] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[762] = {5'd1, 4'd2, 4'd4, 16'd1623};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1623, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[763] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[764] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[765] = {5'd1, 4'd2, 4'd4, 16'd1624};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1624, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[766] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[767] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[768] = {5'd1, 4'd2, 4'd4, 16'd1625};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1625, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[769] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[770] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[771] = {5'd1, 4'd2, 4'd4, 16'd1626};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1626, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[772] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[773] = {5'd0, 4'd8, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 60, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[774] = {5'd1, 4'd2, 4'd4, 16'd1627};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1627, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[775] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[776] = {5'd0, 4'd8, 4'd0, 16'd47};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 47, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[777] = {5'd1, 4'd2, 4'd4, 16'd1628};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1628, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[778] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[779] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[780] = {5'd1, 4'd2, 4'd4, 16'd1629};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1629, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[781] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[782] = {5'd0, 4'd8, 4'd0, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 62, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[783] = {5'd1, 4'd2, 4'd4, 16'd1630};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1630, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[784] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[785] = {5'd0, 4'd8, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 60, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[786] = {5'd1, 4'd2, 4'd4, 16'd1631};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1631, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[787] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[788] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[789] = {5'd1, 4'd2, 4'd4, 16'd1632};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1632, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[790] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[791] = {5'd0, 4'd8, 4'd0, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 62, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[792] = {5'd1, 4'd2, 4'd4, 16'd1633};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1633, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[793] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[794] = {5'd0, 4'd8, 4'd0, 16'd66};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 66, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[795] = {5'd1, 4'd2, 4'd4, 16'd1634};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1634, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[796] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[797] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[798] = {5'd1, 4'd2, 4'd4, 16'd1635};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1635, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[799] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[800] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[801] = {5'd1, 4'd2, 4'd4, 16'd1636};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1636, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[802] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[803] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[804] = {5'd1, 4'd2, 4'd4, 16'd1637};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1637, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[805] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[806] = {5'd0, 4'd8, 4'd0, 16'd111};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 111, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[807] = {5'd1, 4'd2, 4'd4, 16'd1638};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1638, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[808] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[809] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[810] = {5'd1, 4'd2, 4'd4, 16'd1639};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1639, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[811] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[812] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[813] = {5'd1, 4'd2, 4'd4, 16'd1640};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1640, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[814] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[815] = {5'd0, 4'd8, 4'd0, 16'd83};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 83, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[816] = {5'd1, 4'd2, 4'd4, 16'd1641};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1641, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[817] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[818] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[819] = {5'd1, 4'd2, 4'd4, 16'd1642};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1642, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[820] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[821] = {5'd0, 4'd8, 4'd0, 16'd97};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 97, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[822] = {5'd1, 4'd2, 4'd4, 16'd1643};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1643, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[823] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[824] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[825] = {5'd1, 4'd2, 4'd4, 16'd1644};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1644, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[826] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[827] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[828] = {5'd1, 4'd2, 4'd4, 16'd1645};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1645, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[829] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[830] = {5'd0, 4'd8, 4'd0, 16'd115};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 115, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[831] = {5'd1, 4'd2, 4'd4, 16'd1646};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1646, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[832] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[833] = {5'd0, 4'd8, 4'd0, 16'd58};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 58, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[834] = {5'd1, 4'd2, 4'd4, 16'd1647};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1647, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[835] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[836] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[837] = {5'd1, 4'd2, 4'd4, 16'd1648};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1648, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[838] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[839] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[840] = {5'd1, 4'd2, 4'd4, 16'd1649};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1649, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[841] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[842] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[843] = {5'd1, 4'd2, 4'd4, 16'd1650};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1650, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[844] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[845] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[846] = {5'd1, 4'd2, 4'd4, 16'd1651};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1651, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[847] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[848] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[849] = {5'd1, 4'd2, 4'd4, 16'd1652};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1652, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[850] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[851] = {5'd0, 4'd8, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 60, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[852] = {5'd1, 4'd2, 4'd4, 16'd1653};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1653, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[853] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[854] = {5'd0, 4'd8, 4'd0, 16'd47};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 47, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[855] = {5'd1, 4'd2, 4'd4, 16'd1654};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1654, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[856] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[857] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[858] = {5'd1, 4'd2, 4'd4, 16'd1655};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1655, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[859] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[860] = {5'd0, 4'd8, 4'd0, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 62, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[861] = {5'd1, 4'd2, 4'd4, 16'd1656};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1656, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[862] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[863] = {5'd0, 4'd8, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 60, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[864] = {5'd1, 4'd2, 4'd4, 16'd1657};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1657, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[865] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[866] = {5'd0, 4'd8, 4'd0, 16'd102};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 102, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[867] = {5'd1, 4'd2, 4'd4, 16'd1658};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1658, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[868] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[869] = {5'd0, 4'd8, 4'd0, 16'd111};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 111, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[870] = {5'd1, 4'd2, 4'd4, 16'd1659};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1659, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[871] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[872] = {5'd0, 4'd8, 4'd0, 16'd114};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 114, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[873] = {5'd1, 4'd2, 4'd4, 16'd1660};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1660, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[874] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[875] = {5'd0, 4'd8, 4'd0, 16'd109};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 109, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[876] = {5'd1, 4'd2, 4'd4, 16'd1661};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1661, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[877] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[878] = {5'd0, 4'd8, 4'd0, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 62, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[879] = {5'd1, 4'd2, 4'd4, 16'd1662};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1662, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[880] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[881] = {5'd0, 4'd8, 4'd0, 16'd9};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 9, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[882] = {5'd1, 4'd2, 4'd4, 16'd1663};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1663, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[883] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[884] = {5'd0, 4'd8, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 60, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[885] = {5'd1, 4'd2, 4'd4, 16'd1664};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1664, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[886] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[887] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[888] = {5'd1, 4'd2, 4'd4, 16'd1665};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1665, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[889] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[890] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[891] = {5'd1, 4'd2, 4'd4, 16'd1666};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1666, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[892] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[893] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[894] = {5'd1, 4'd2, 4'd4, 16'd1667};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1667, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[895] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[896] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[897] = {5'd1, 4'd2, 4'd4, 16'd1668};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1668, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[898] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[899] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[900] = {5'd1, 4'd2, 4'd4, 16'd1669};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1669, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[901] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[902] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[903] = {5'd1, 4'd2, 4'd4, 16'd1670};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1670, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[904] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[905] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[906] = {5'd1, 4'd2, 4'd4, 16'd1671};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1671, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[907] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[908] = {5'd0, 4'd8, 4'd0, 16'd121};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 121, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[909] = {5'd1, 4'd2, 4'd4, 16'd1672};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1672, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[910] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[911] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[912] = {5'd1, 4'd2, 4'd4, 16'd1673};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1673, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[913] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[914] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[915] = {5'd1, 4'd2, 4'd4, 16'd1674};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1674, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[916] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[917] = {5'd0, 4'd8, 4'd0, 16'd61};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 61, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[918] = {5'd1, 4'd2, 4'd4, 16'd1675};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1675, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[919] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[920] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[921] = {5'd1, 4'd2, 4'd4, 16'd1676};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1676, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[922] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[923] = {5'd0, 4'd8, 4'd0, 16'd99};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 99, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[924] = {5'd1, 4'd2, 4'd4, 16'd1677};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1677, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[925] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[926] = {5'd0, 4'd8, 4'd0, 16'd104};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 104, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[927] = {5'd1, 4'd2, 4'd4, 16'd1678};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1678, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[928] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[929] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[930] = {5'd1, 4'd2, 4'd4, 16'd1679};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1679, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[931] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[932] = {5'd0, 4'd8, 4'd0, 16'd99};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 99, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[933] = {5'd1, 4'd2, 4'd4, 16'd1680};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1680, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[934] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[935] = {5'd0, 4'd8, 4'd0, 16'd107};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 107, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[936] = {5'd1, 4'd2, 4'd4, 16'd1681};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1681, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[937] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[938] = {5'd0, 4'd8, 4'd0, 16'd98};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 98, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[939] = {5'd1, 4'd2, 4'd4, 16'd1682};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1682, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[940] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[941] = {5'd0, 4'd8, 4'd0, 16'd111};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 111, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[942] = {5'd1, 4'd2, 4'd4, 16'd1683};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1683, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[943] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[944] = {5'd0, 4'd8, 4'd0, 16'd120};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 120, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[945] = {5'd1, 4'd2, 4'd4, 16'd1684};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1684, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[946] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[947] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[948] = {5'd1, 4'd2, 4'd4, 16'd1685};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1685, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[949] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[950] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[951] = {5'd1, 4'd2, 4'd4, 16'd1686};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1686, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[952] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[953] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[954] = {5'd1, 4'd2, 4'd4, 16'd1687};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1687, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[955] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[956] = {5'd0, 4'd8, 4'd0, 16'd97};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 97, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[957] = {5'd1, 4'd2, 4'd4, 16'd1688};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1688, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[958] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[959] = {5'd0, 4'd8, 4'd0, 16'd109};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 109, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[960] = {5'd1, 4'd2, 4'd4, 16'd1689};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1689, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[961] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[962] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[963] = {5'd1, 4'd2, 4'd4, 16'd1690};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1690, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[964] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[965] = {5'd0, 4'd8, 4'd0, 16'd61};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 61, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[966] = {5'd1, 4'd2, 4'd4, 16'd1691};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1691, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[967] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[968] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[969] = {5'd1, 4'd2, 4'd4, 16'd1692};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1692, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[970] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[971] = {5'd0, 4'd8, 4'd0, 16'd108};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 108, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[972] = {5'd1, 4'd2, 4'd4, 16'd1693};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1693, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[973] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[974] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[975] = {5'd1, 4'd2, 4'd4, 16'd1694};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1694, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[976] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[977] = {5'd0, 4'd8, 4'd0, 16'd100};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 100, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[978] = {5'd1, 4'd2, 4'd4, 16'd1695};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1695, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[979] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[980] = {5'd0, 4'd8, 4'd0, 16'd49};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 49, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[981] = {5'd1, 4'd2, 4'd4, 16'd1696};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1696, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[982] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[983] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[984] = {5'd1, 4'd2, 4'd4, 16'd1697};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1697, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[985] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[986] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[987] = {5'd1, 4'd2, 4'd4, 16'd1698};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1698, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[988] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[989] = {5'd0, 4'd8, 4'd0, 16'd118};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 118, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[990] = {5'd1, 4'd2, 4'd4, 16'd1699};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1699, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[991] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[992] = {5'd0, 4'd8, 4'd0, 16'd97};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 97, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[993] = {5'd1, 4'd2, 4'd4, 16'd1700};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1700, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[994] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[995] = {5'd0, 4'd8, 4'd0, 16'd108};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 108, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[996] = {5'd1, 4'd2, 4'd4, 16'd1701};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1701, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[997] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[998] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[999] = {5'd1, 4'd2, 4'd4, 16'd1702};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1702, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1000] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1001] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1002] = {5'd1, 4'd2, 4'd4, 16'd1703};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1703, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1003] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1004] = {5'd0, 4'd8, 4'd0, 16'd61};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 61, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1005] = {5'd1, 4'd2, 4'd4, 16'd1704};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1704, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1006] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1007] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1008] = {5'd1, 4'd2, 4'd4, 16'd1705};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1705, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1009] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1010] = {5'd0, 4'd8, 4'd0, 16'd65};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 65, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1011] = {5'd1, 4'd2, 4'd4, 16'd1706};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1706, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1012] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1013] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1014] = {5'd1, 4'd2, 4'd4, 16'd1707};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1707, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1015] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1016] = {5'd0, 4'd8, 4'd0, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 62, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1017] = {5'd1, 4'd2, 4'd4, 16'd1708};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1708, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1018] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1019] = {5'd0, 4'd8, 4'd0, 16'd108};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 108, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1020] = {5'd1, 4'd2, 4'd4, 16'd1709};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1709, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1021] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1022] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1023] = {5'd1, 4'd2, 4'd4, 16'd1710};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1710, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1024] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1025] = {5'd0, 4'd8, 4'd0, 16'd100};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 100, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1026] = {5'd1, 4'd2, 4'd4, 16'd1711};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1711, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1027] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1028] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1029] = {5'd1, 4'd2, 4'd4, 16'd1712};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1712, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1030] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1031] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1032] = {5'd1, 4'd2, 4'd4, 16'd1713};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1713, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1033] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1034] = {5'd0, 4'd8, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 60, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1035] = {5'd1, 4'd2, 4'd4, 16'd1714};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1714, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1036] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1037] = {5'd0, 4'd8, 4'd0, 16'd47};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 47, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1038] = {5'd1, 4'd2, 4'd4, 16'd1715};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1715, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1039] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1040] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1041] = {5'd1, 4'd2, 4'd4, 16'd1716};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1716, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1042] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1043] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1044] = {5'd1, 4'd2, 4'd4, 16'd1717};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1717, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1045] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1046] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1047] = {5'd1, 4'd2, 4'd4, 16'd1718};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1718, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1048] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1049] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1050] = {5'd1, 4'd2, 4'd4, 16'd1719};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1719, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1051] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1052] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1053] = {5'd1, 4'd2, 4'd4, 16'd1720};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1720, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1054] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1055] = {5'd0, 4'd8, 4'd0, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 62, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1056] = {5'd1, 4'd2, 4'd4, 16'd1721};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1721, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1057] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1058] = {5'd0, 4'd8, 4'd0, 16'd9};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 9, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1059] = {5'd1, 4'd2, 4'd4, 16'd1722};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1722, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1060] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1061] = {5'd0, 4'd8, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 60, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1062] = {5'd1, 4'd2, 4'd4, 16'd1723};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1723, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1063] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1064] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1065] = {5'd1, 4'd2, 4'd4, 16'd1724};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1724, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1066] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1067] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1068] = {5'd1, 4'd2, 4'd4, 16'd1725};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1725, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1069] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1070] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1071] = {5'd1, 4'd2, 4'd4, 16'd1726};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1726, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1072] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1073] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1074] = {5'd1, 4'd2, 4'd4, 16'd1727};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1727, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1075] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1076] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1077] = {5'd1, 4'd2, 4'd4, 16'd1728};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1728, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1078] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1079] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1080] = {5'd1, 4'd2, 4'd4, 16'd1729};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1729, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1081] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1082] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1083] = {5'd1, 4'd2, 4'd4, 16'd1730};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1730, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1084] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1085] = {5'd0, 4'd8, 4'd0, 16'd121};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 121, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1086] = {5'd1, 4'd2, 4'd4, 16'd1731};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1731, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1087] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1088] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1089] = {5'd1, 4'd2, 4'd4, 16'd1732};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1732, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1090] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1091] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1092] = {5'd1, 4'd2, 4'd4, 16'd1733};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1733, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1093] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1094] = {5'd0, 4'd8, 4'd0, 16'd61};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 61, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1095] = {5'd1, 4'd2, 4'd4, 16'd1734};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1734, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1096] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1097] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1098] = {5'd1, 4'd2, 4'd4, 16'd1735};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1735, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1099] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1100] = {5'd0, 4'd8, 4'd0, 16'd99};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 99, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1101] = {5'd1, 4'd2, 4'd4, 16'd1736};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1736, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1102] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1103] = {5'd0, 4'd8, 4'd0, 16'd104};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 104, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1104] = {5'd1, 4'd2, 4'd4, 16'd1737};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1737, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1105] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1106] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1107] = {5'd1, 4'd2, 4'd4, 16'd1738};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1738, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1108] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1109] = {5'd0, 4'd8, 4'd0, 16'd99};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 99, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1110] = {5'd1, 4'd2, 4'd4, 16'd1739};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1739, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1111] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1112] = {5'd0, 4'd8, 4'd0, 16'd107};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 107, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1113] = {5'd1, 4'd2, 4'd4, 16'd1740};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1740, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1114] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1115] = {5'd0, 4'd8, 4'd0, 16'd98};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 98, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1116] = {5'd1, 4'd2, 4'd4, 16'd1741};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1741, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1117] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1118] = {5'd0, 4'd8, 4'd0, 16'd111};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 111, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1119] = {5'd1, 4'd2, 4'd4, 16'd1742};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1742, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1120] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1121] = {5'd0, 4'd8, 4'd0, 16'd120};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 120, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1122] = {5'd1, 4'd2, 4'd4, 16'd1743};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1743, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1123] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1124] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1125] = {5'd1, 4'd2, 4'd4, 16'd1744};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1744, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1126] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1127] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1128] = {5'd1, 4'd2, 4'd4, 16'd1745};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1745, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1129] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1130] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1131] = {5'd1, 4'd2, 4'd4, 16'd1746};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1746, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1132] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1133] = {5'd0, 4'd8, 4'd0, 16'd97};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 97, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1134] = {5'd1, 4'd2, 4'd4, 16'd1747};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1747, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1135] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1136] = {5'd0, 4'd8, 4'd0, 16'd109};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 109, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1137] = {5'd1, 4'd2, 4'd4, 16'd1748};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1748, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1138] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1139] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1140] = {5'd1, 4'd2, 4'd4, 16'd1749};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1749, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1141] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1142] = {5'd0, 4'd8, 4'd0, 16'd61};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 61, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1143] = {5'd1, 4'd2, 4'd4, 16'd1750};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1750, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1144] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1145] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1146] = {5'd1, 4'd2, 4'd4, 16'd1751};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1751, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1147] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1148] = {5'd0, 4'd8, 4'd0, 16'd108};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 108, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1149] = {5'd1, 4'd2, 4'd4, 16'd1752};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1752, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1150] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1151] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1152] = {5'd1, 4'd2, 4'd4, 16'd1753};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1753, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1153] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1154] = {5'd0, 4'd8, 4'd0, 16'd100};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 100, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1155] = {5'd1, 4'd2, 4'd4, 16'd1754};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1754, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1156] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1157] = {5'd0, 4'd8, 4'd0, 16'd50};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 50, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1158] = {5'd1, 4'd2, 4'd4, 16'd1755};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1755, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1159] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1160] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1161] = {5'd1, 4'd2, 4'd4, 16'd1756};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1756, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1162] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1163] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1164] = {5'd1, 4'd2, 4'd4, 16'd1757};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1757, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1165] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1166] = {5'd0, 4'd8, 4'd0, 16'd118};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 118, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1167] = {5'd1, 4'd2, 4'd4, 16'd1758};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1758, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1168] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1169] = {5'd0, 4'd8, 4'd0, 16'd97};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 97, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1170] = {5'd1, 4'd2, 4'd4, 16'd1759};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1759, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1171] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1172] = {5'd0, 4'd8, 4'd0, 16'd108};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 108, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1173] = {5'd1, 4'd2, 4'd4, 16'd1760};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1760, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1174] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1175] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1176] = {5'd1, 4'd2, 4'd4, 16'd1761};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1761, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1177] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1178] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1179] = {5'd1, 4'd2, 4'd4, 16'd1762};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1762, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1180] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1181] = {5'd0, 4'd8, 4'd0, 16'd61};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 61, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1182] = {5'd1, 4'd2, 4'd4, 16'd1763};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1763, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1183] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1184] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1185] = {5'd1, 4'd2, 4'd4, 16'd1764};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1764, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1186] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1187] = {5'd0, 4'd8, 4'd0, 16'd66};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 66, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1188] = {5'd1, 4'd2, 4'd4, 16'd1765};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1765, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1189] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1190] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1191] = {5'd1, 4'd2, 4'd4, 16'd1766};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1766, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1192] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1193] = {5'd0, 4'd8, 4'd0, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 62, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1194] = {5'd1, 4'd2, 4'd4, 16'd1767};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1767, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1195] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1196] = {5'd0, 4'd8, 4'd0, 16'd108};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 108, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1197] = {5'd1, 4'd2, 4'd4, 16'd1768};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1768, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1198] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1199] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1200] = {5'd1, 4'd2, 4'd4, 16'd1769};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1769, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1201] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1202] = {5'd0, 4'd8, 4'd0, 16'd100};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 100, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1203] = {5'd1, 4'd2, 4'd4, 16'd1770};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1770, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1204] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1205] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1206] = {5'd1, 4'd2, 4'd4, 16'd1771};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1771, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1207] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1208] = {5'd0, 4'd8, 4'd0, 16'd49};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 49, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1209] = {5'd1, 4'd2, 4'd4, 16'd1772};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1772, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1210] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1211] = {5'd0, 4'd8, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 60, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1212] = {5'd1, 4'd2, 4'd4, 16'd1773};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1773, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1213] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1214] = {5'd0, 4'd8, 4'd0, 16'd47};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 47, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1215] = {5'd1, 4'd2, 4'd4, 16'd1774};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1774, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1216] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1217] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1218] = {5'd1, 4'd2, 4'd4, 16'd1775};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1775, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1219] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1220] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1221] = {5'd1, 4'd2, 4'd4, 16'd1776};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1776, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1222] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1223] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1224] = {5'd1, 4'd2, 4'd4, 16'd1777};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1777, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1225] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1226] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1227] = {5'd1, 4'd2, 4'd4, 16'd1778};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1778, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1228] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1229] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1230] = {5'd1, 4'd2, 4'd4, 16'd1779};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1779, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1231] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1232] = {5'd0, 4'd8, 4'd0, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 62, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1233] = {5'd1, 4'd2, 4'd4, 16'd1780};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1780, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1234] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1235] = {5'd0, 4'd8, 4'd0, 16'd9};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 9, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1236] = {5'd1, 4'd2, 4'd4, 16'd1781};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1781, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1237] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1238] = {5'd0, 4'd8, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 60, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1239] = {5'd1, 4'd2, 4'd4, 16'd1782};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1782, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1240] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1241] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1242] = {5'd1, 4'd2, 4'd4, 16'd1783};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1783, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1243] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1244] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1245] = {5'd1, 4'd2, 4'd4, 16'd1784};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1784, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1246] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1247] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1248] = {5'd1, 4'd2, 4'd4, 16'd1785};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1785, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1249] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1250] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1251] = {5'd1, 4'd2, 4'd4, 16'd1786};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1786, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1252] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1253] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1254] = {5'd1, 4'd2, 4'd4, 16'd1787};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1787, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1255] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1256] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1257] = {5'd1, 4'd2, 4'd4, 16'd1788};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1788, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1258] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1259] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1260] = {5'd1, 4'd2, 4'd4, 16'd1789};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1789, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1261] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1262] = {5'd0, 4'd8, 4'd0, 16'd121};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 121, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1263] = {5'd1, 4'd2, 4'd4, 16'd1790};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1790, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1264] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1265] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1266] = {5'd1, 4'd2, 4'd4, 16'd1791};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1791, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1267] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1268] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1269] = {5'd1, 4'd2, 4'd4, 16'd1792};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1792, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1270] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1271] = {5'd0, 4'd8, 4'd0, 16'd61};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 61, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1272] = {5'd1, 4'd2, 4'd4, 16'd1793};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1793, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1273] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1274] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1275] = {5'd1, 4'd2, 4'd4, 16'd1794};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1794, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1276] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1277] = {5'd0, 4'd8, 4'd0, 16'd99};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 99, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1278] = {5'd1, 4'd2, 4'd4, 16'd1795};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1795, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1279] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1280] = {5'd0, 4'd8, 4'd0, 16'd104};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 104, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1281] = {5'd1, 4'd2, 4'd4, 16'd1796};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1796, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1282] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1283] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1284] = {5'd1, 4'd2, 4'd4, 16'd1797};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1797, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1285] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1286] = {5'd0, 4'd8, 4'd0, 16'd99};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 99, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1287] = {5'd1, 4'd2, 4'd4, 16'd1798};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1798, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1288] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1289] = {5'd0, 4'd8, 4'd0, 16'd107};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 107, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1290] = {5'd1, 4'd2, 4'd4, 16'd1799};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1799, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1291] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1292] = {5'd0, 4'd8, 4'd0, 16'd98};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 98, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1293] = {5'd1, 4'd2, 4'd4, 16'd1800};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1800, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1294] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1295] = {5'd0, 4'd8, 4'd0, 16'd111};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 111, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1296] = {5'd1, 4'd2, 4'd4, 16'd1801};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1801, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1297] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1298] = {5'd0, 4'd8, 4'd0, 16'd120};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 120, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1299] = {5'd1, 4'd2, 4'd4, 16'd1802};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1802, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1300] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1301] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1302] = {5'd1, 4'd2, 4'd4, 16'd1803};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1803, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1303] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1304] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1305] = {5'd1, 4'd2, 4'd4, 16'd1804};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1804, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1306] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1307] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1308] = {5'd1, 4'd2, 4'd4, 16'd1805};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1805, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1309] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1310] = {5'd0, 4'd8, 4'd0, 16'd97};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 97, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1311] = {5'd1, 4'd2, 4'd4, 16'd1806};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1806, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1312] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1313] = {5'd0, 4'd8, 4'd0, 16'd109};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 109, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1314] = {5'd1, 4'd2, 4'd4, 16'd1807};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1807, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1315] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1316] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1317] = {5'd1, 4'd2, 4'd4, 16'd1808};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1808, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1318] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1319] = {5'd0, 4'd8, 4'd0, 16'd61};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 61, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1320] = {5'd1, 4'd2, 4'd4, 16'd1809};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1809, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1321] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1322] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1323] = {5'd1, 4'd2, 4'd4, 16'd1810};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1810, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1324] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1325] = {5'd0, 4'd8, 4'd0, 16'd108};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 108, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1326] = {5'd1, 4'd2, 4'd4, 16'd1811};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1811, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1327] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1328] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1329] = {5'd1, 4'd2, 4'd4, 16'd1812};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1812, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1330] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1331] = {5'd0, 4'd8, 4'd0, 16'd100};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 100, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1332] = {5'd1, 4'd2, 4'd4, 16'd1813};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1813, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1333] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1334] = {5'd0, 4'd8, 4'd0, 16'd51};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 51, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1335] = {5'd1, 4'd2, 4'd4, 16'd1814};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1814, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1336] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1337] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1338] = {5'd1, 4'd2, 4'd4, 16'd1815};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1815, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1339] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1340] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1341] = {5'd1, 4'd2, 4'd4, 16'd1816};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1816, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1342] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1343] = {5'd0, 4'd8, 4'd0, 16'd118};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 118, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1344] = {5'd1, 4'd2, 4'd4, 16'd1817};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1817, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1345] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1346] = {5'd0, 4'd8, 4'd0, 16'd97};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 97, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1347] = {5'd1, 4'd2, 4'd4, 16'd1818};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1818, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1348] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1349] = {5'd0, 4'd8, 4'd0, 16'd108};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 108, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1350] = {5'd1, 4'd2, 4'd4, 16'd1819};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1819, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1351] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1352] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1353] = {5'd1, 4'd2, 4'd4, 16'd1820};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1820, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1354] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1355] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1356] = {5'd1, 4'd2, 4'd4, 16'd1821};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1821, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1357] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1358] = {5'd0, 4'd8, 4'd0, 16'd61};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 61, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1359] = {5'd1, 4'd2, 4'd4, 16'd1822};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1822, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1360] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1361] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1362] = {5'd1, 4'd2, 4'd4, 16'd1823};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1823, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1363] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1364] = {5'd0, 4'd8, 4'd0, 16'd67};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 67, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1365] = {5'd1, 4'd2, 4'd4, 16'd1824};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1824, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1366] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1367] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1368] = {5'd1, 4'd2, 4'd4, 16'd1825};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1825, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1369] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1370] = {5'd0, 4'd8, 4'd0, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 62, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1371] = {5'd1, 4'd2, 4'd4, 16'd1826};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1826, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1372] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1373] = {5'd0, 4'd8, 4'd0, 16'd108};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 108, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1374] = {5'd1, 4'd2, 4'd4, 16'd1827};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1827, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1375] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1376] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1377] = {5'd1, 4'd2, 4'd4, 16'd1828};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1828, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1378] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1379] = {5'd0, 4'd8, 4'd0, 16'd100};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 100, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1380] = {5'd1, 4'd2, 4'd4, 16'd1829};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1829, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1381] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1382] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1383] = {5'd1, 4'd2, 4'd4, 16'd1830};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1830, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1384] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1385] = {5'd0, 4'd8, 4'd0, 16'd50};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 50, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1386] = {5'd1, 4'd2, 4'd4, 16'd1831};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1831, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1387] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1388] = {5'd0, 4'd8, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 60, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1389] = {5'd1, 4'd2, 4'd4, 16'd1832};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1832, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1390] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1391] = {5'd0, 4'd8, 4'd0, 16'd47};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 47, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1392] = {5'd1, 4'd2, 4'd4, 16'd1833};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1833, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1393] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1394] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1395] = {5'd1, 4'd2, 4'd4, 16'd1834};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1834, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1396] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1397] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1398] = {5'd1, 4'd2, 4'd4, 16'd1835};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1835, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1399] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1400] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1401] = {5'd1, 4'd2, 4'd4, 16'd1836};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1836, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1402] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1403] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1404] = {5'd1, 4'd2, 4'd4, 16'd1837};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1837, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1405] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1406] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1407] = {5'd1, 4'd2, 4'd4, 16'd1838};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1838, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1408] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1409] = {5'd0, 4'd8, 4'd0, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 62, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1410] = {5'd1, 4'd2, 4'd4, 16'd1839};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1839, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1411] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1412] = {5'd0, 4'd8, 4'd0, 16'd9};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 9, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1413] = {5'd1, 4'd2, 4'd4, 16'd1840};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1840, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1414] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1415] = {5'd0, 4'd8, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 60, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1416] = {5'd1, 4'd2, 4'd4, 16'd1841};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1841, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1417] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1418] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1419] = {5'd1, 4'd2, 4'd4, 16'd1842};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1842, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1420] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1421] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1422] = {5'd1, 4'd2, 4'd4, 16'd1843};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1843, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1423] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1424] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1425] = {5'd1, 4'd2, 4'd4, 16'd1844};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1844, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1426] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1427] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1428] = {5'd1, 4'd2, 4'd4, 16'd1845};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1845, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1429] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1430] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1431] = {5'd1, 4'd2, 4'd4, 16'd1846};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1846, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1432] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1433] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1434] = {5'd1, 4'd2, 4'd4, 16'd1847};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1847, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1435] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1436] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1437] = {5'd1, 4'd2, 4'd4, 16'd1848};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1848, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1438] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1439] = {5'd0, 4'd8, 4'd0, 16'd121};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 121, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1440] = {5'd1, 4'd2, 4'd4, 16'd1849};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1849, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1441] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1442] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1443] = {5'd1, 4'd2, 4'd4, 16'd1850};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1850, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1444] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1445] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1446] = {5'd1, 4'd2, 4'd4, 16'd1851};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1851, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1447] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1448] = {5'd0, 4'd8, 4'd0, 16'd61};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 61, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1449] = {5'd1, 4'd2, 4'd4, 16'd1852};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1852, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1450] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1451] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1452] = {5'd1, 4'd2, 4'd4, 16'd1853};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1853, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1453] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1454] = {5'd0, 4'd8, 4'd0, 16'd99};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 99, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1455] = {5'd1, 4'd2, 4'd4, 16'd1854};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1854, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1456] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1457] = {5'd0, 4'd8, 4'd0, 16'd104};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 104, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1458] = {5'd1, 4'd2, 4'd4, 16'd1855};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1855, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1459] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1460] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1461] = {5'd1, 4'd2, 4'd4, 16'd1856};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1856, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1462] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1463] = {5'd0, 4'd8, 4'd0, 16'd99};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 99, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1464] = {5'd1, 4'd2, 4'd4, 16'd1857};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1857, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1465] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1466] = {5'd0, 4'd8, 4'd0, 16'd107};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 107, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1467] = {5'd1, 4'd2, 4'd4, 16'd1858};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1858, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1468] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1469] = {5'd0, 4'd8, 4'd0, 16'd98};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 98, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1470] = {5'd1, 4'd2, 4'd4, 16'd1859};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1859, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1471] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1472] = {5'd0, 4'd8, 4'd0, 16'd111};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 111, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1473] = {5'd1, 4'd2, 4'd4, 16'd1860};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1860, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1474] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1475] = {5'd0, 4'd8, 4'd0, 16'd120};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 120, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1476] = {5'd1, 4'd2, 4'd4, 16'd1861};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1861, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1477] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1478] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1479] = {5'd1, 4'd2, 4'd4, 16'd1862};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1862, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1480] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1481] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1482] = {5'd1, 4'd2, 4'd4, 16'd1863};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1863, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1483] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1484] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1485] = {5'd1, 4'd2, 4'd4, 16'd1864};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1864, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1486] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1487] = {5'd0, 4'd8, 4'd0, 16'd97};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 97, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1488] = {5'd1, 4'd2, 4'd4, 16'd1865};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1865, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1489] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1490] = {5'd0, 4'd8, 4'd0, 16'd109};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 109, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1491] = {5'd1, 4'd2, 4'd4, 16'd1866};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1866, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1492] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1493] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1494] = {5'd1, 4'd2, 4'd4, 16'd1867};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1867, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1495] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1496] = {5'd0, 4'd8, 4'd0, 16'd61};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 61, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1497] = {5'd1, 4'd2, 4'd4, 16'd1868};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1868, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1498] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1499] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1500] = {5'd1, 4'd2, 4'd4, 16'd1869};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1869, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1501] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1502] = {5'd0, 4'd8, 4'd0, 16'd108};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 108, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1503] = {5'd1, 4'd2, 4'd4, 16'd1870};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1870, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1504] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1505] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1506] = {5'd1, 4'd2, 4'd4, 16'd1871};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1871, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1507] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1508] = {5'd0, 4'd8, 4'd0, 16'd100};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 100, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1509] = {5'd1, 4'd2, 4'd4, 16'd1872};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1872, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1510] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1511] = {5'd0, 4'd8, 4'd0, 16'd52};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 52, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1512] = {5'd1, 4'd2, 4'd4, 16'd1873};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1873, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1513] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1514] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1515] = {5'd1, 4'd2, 4'd4, 16'd1874};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1874, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1516] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1517] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1518] = {5'd1, 4'd2, 4'd4, 16'd1875};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1875, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1519] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1520] = {5'd0, 4'd8, 4'd0, 16'd118};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 118, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1521] = {5'd1, 4'd2, 4'd4, 16'd1876};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1876, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1522] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1523] = {5'd0, 4'd8, 4'd0, 16'd97};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 97, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1524] = {5'd1, 4'd2, 4'd4, 16'd1877};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1877, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1525] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1526] = {5'd0, 4'd8, 4'd0, 16'd108};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 108, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1527] = {5'd1, 4'd2, 4'd4, 16'd1878};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1878, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1528] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1529] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1530] = {5'd1, 4'd2, 4'd4, 16'd1879};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1879, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1531] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1532] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1533] = {5'd1, 4'd2, 4'd4, 16'd1880};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1880, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1534] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1535] = {5'd0, 4'd8, 4'd0, 16'd61};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 61, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1536] = {5'd1, 4'd2, 4'd4, 16'd1881};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1881, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1537] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1538] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1539] = {5'd1, 4'd2, 4'd4, 16'd1882};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1882, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1540] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1541] = {5'd0, 4'd8, 4'd0, 16'd68};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 68, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1542] = {5'd1, 4'd2, 4'd4, 16'd1883};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1883, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1543] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1544] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1545] = {5'd1, 4'd2, 4'd4, 16'd1884};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1884, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1546] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1547] = {5'd0, 4'd8, 4'd0, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 62, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1548] = {5'd1, 4'd2, 4'd4, 16'd1885};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1885, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1549] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1550] = {5'd0, 4'd8, 4'd0, 16'd108};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 108, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1551] = {5'd1, 4'd2, 4'd4, 16'd1886};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1886, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1552] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1553] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1554] = {5'd1, 4'd2, 4'd4, 16'd1887};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1887, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1555] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1556] = {5'd0, 4'd8, 4'd0, 16'd100};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 100, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1557] = {5'd1, 4'd2, 4'd4, 16'd1888};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1888, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1558] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1559] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1560] = {5'd1, 4'd2, 4'd4, 16'd1889};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1889, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1561] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1562] = {5'd0, 4'd8, 4'd0, 16'd51};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 51, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1563] = {5'd1, 4'd2, 4'd4, 16'd1890};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1890, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1564] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1565] = {5'd0, 4'd8, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 60, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1566] = {5'd1, 4'd2, 4'd4, 16'd1891};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1891, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1567] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1568] = {5'd0, 4'd8, 4'd0, 16'd47};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 47, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1569] = {5'd1, 4'd2, 4'd4, 16'd1892};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1892, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1570] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1571] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1572] = {5'd1, 4'd2, 4'd4, 16'd1893};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1893, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1573] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1574] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1575] = {5'd1, 4'd2, 4'd4, 16'd1894};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1894, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1576] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1577] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1578] = {5'd1, 4'd2, 4'd4, 16'd1895};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1895, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1579] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1580] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1581] = {5'd1, 4'd2, 4'd4, 16'd1896};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1896, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1582] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1583] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1584] = {5'd1, 4'd2, 4'd4, 16'd1897};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1897, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1585] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1586] = {5'd0, 4'd8, 4'd0, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 62, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1587] = {5'd1, 4'd2, 4'd4, 16'd1898};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1898, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1588] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1589] = {5'd0, 4'd8, 4'd0, 16'd9};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 9, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1590] = {5'd1, 4'd2, 4'd4, 16'd1899};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1899, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1591] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1592] = {5'd0, 4'd8, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 60, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1593] = {5'd1, 4'd2, 4'd4, 16'd1900};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1900, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1594] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1595] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1596] = {5'd1, 4'd2, 4'd4, 16'd1901};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1901, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1597] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1598] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1599] = {5'd1, 4'd2, 4'd4, 16'd1902};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1902, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1600] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1601] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1602] = {5'd1, 4'd2, 4'd4, 16'd1903};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1903, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1603] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1604] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1605] = {5'd1, 4'd2, 4'd4, 16'd1904};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1904, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1606] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1607] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1608] = {5'd1, 4'd2, 4'd4, 16'd1905};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1905, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1609] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1610] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1611] = {5'd1, 4'd2, 4'd4, 16'd1906};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1906, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1612] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1613] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1614] = {5'd1, 4'd2, 4'd4, 16'd1907};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1907, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1615] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1616] = {5'd0, 4'd8, 4'd0, 16'd121};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 121, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1617] = {5'd1, 4'd2, 4'd4, 16'd1908};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1908, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1618] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1619] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1620] = {5'd1, 4'd2, 4'd4, 16'd1909};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1909, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1621] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1622] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1623] = {5'd1, 4'd2, 4'd4, 16'd1910};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1910, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1624] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1625] = {5'd0, 4'd8, 4'd0, 16'd61};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 61, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1626] = {5'd1, 4'd2, 4'd4, 16'd1911};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1911, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1627] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1628] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1629] = {5'd1, 4'd2, 4'd4, 16'd1912};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1912, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1630] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1631] = {5'd0, 4'd8, 4'd0, 16'd99};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 99, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1632] = {5'd1, 4'd2, 4'd4, 16'd1913};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1913, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1633] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1634] = {5'd0, 4'd8, 4'd0, 16'd104};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 104, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1635] = {5'd1, 4'd2, 4'd4, 16'd1914};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1914, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1636] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1637] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1638] = {5'd1, 4'd2, 4'd4, 16'd1915};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1915, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1639] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1640] = {5'd0, 4'd8, 4'd0, 16'd99};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 99, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1641] = {5'd1, 4'd2, 4'd4, 16'd1916};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1916, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1642] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1643] = {5'd0, 4'd8, 4'd0, 16'd107};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 107, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1644] = {5'd1, 4'd2, 4'd4, 16'd1917};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1917, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1645] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1646] = {5'd0, 4'd8, 4'd0, 16'd98};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 98, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1647] = {5'd1, 4'd2, 4'd4, 16'd1918};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1918, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1648] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1649] = {5'd0, 4'd8, 4'd0, 16'd111};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 111, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1650] = {5'd1, 4'd2, 4'd4, 16'd1919};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1919, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1651] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1652] = {5'd0, 4'd8, 4'd0, 16'd120};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 120, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1653] = {5'd1, 4'd2, 4'd4, 16'd1920};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1920, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1654] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1655] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1656] = {5'd1, 4'd2, 4'd4, 16'd1921};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1921, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1657] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1658] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1659] = {5'd1, 4'd2, 4'd4, 16'd1922};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1922, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1660] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1661] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1662] = {5'd1, 4'd2, 4'd4, 16'd1923};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1923, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1663] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1664] = {5'd0, 4'd8, 4'd0, 16'd97};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 97, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1665] = {5'd1, 4'd2, 4'd4, 16'd1924};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1924, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1666] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1667] = {5'd0, 4'd8, 4'd0, 16'd109};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 109, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1668] = {5'd1, 4'd2, 4'd4, 16'd1925};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1925, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1669] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1670] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1671] = {5'd1, 4'd2, 4'd4, 16'd1926};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1926, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1672] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1673] = {5'd0, 4'd8, 4'd0, 16'd61};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 61, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1674] = {5'd1, 4'd2, 4'd4, 16'd1927};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1927, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1675] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1676] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1677] = {5'd1, 4'd2, 4'd4, 16'd1928};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1928, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1678] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1679] = {5'd0, 4'd8, 4'd0, 16'd108};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 108, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1680] = {5'd1, 4'd2, 4'd4, 16'd1929};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1929, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1681] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1682] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1683] = {5'd1, 4'd2, 4'd4, 16'd1930};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1930, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1684] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1685] = {5'd0, 4'd8, 4'd0, 16'd100};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 100, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1686] = {5'd1, 4'd2, 4'd4, 16'd1931};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1931, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1687] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1688] = {5'd0, 4'd8, 4'd0, 16'd52};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 52, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1689] = {5'd1, 4'd2, 4'd4, 16'd1932};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1932, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1690] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1691] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1692] = {5'd1, 4'd2, 4'd4, 16'd1933};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1933, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1693] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1694] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1695] = {5'd1, 4'd2, 4'd4, 16'd1934};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1934, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1696] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1697] = {5'd0, 4'd8, 4'd0, 16'd118};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 118, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1698] = {5'd1, 4'd2, 4'd4, 16'd1935};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1935, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1699] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1700] = {5'd0, 4'd8, 4'd0, 16'd97};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 97, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1701] = {5'd1, 4'd2, 4'd4, 16'd1936};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1936, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1702] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1703] = {5'd0, 4'd8, 4'd0, 16'd108};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 108, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1704] = {5'd1, 4'd2, 4'd4, 16'd1937};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1937, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1705] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1706] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1707] = {5'd1, 4'd2, 4'd4, 16'd1938};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1938, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1708] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1709] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1710] = {5'd1, 4'd2, 4'd4, 16'd1939};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1939, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1711] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1712] = {5'd0, 4'd8, 4'd0, 16'd61};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 61, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1713] = {5'd1, 4'd2, 4'd4, 16'd1940};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1940, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1714] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1715] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1716] = {5'd1, 4'd2, 4'd4, 16'd1941};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1941, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1717] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1718] = {5'd0, 4'd8, 4'd0, 16'd69};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 69, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1719] = {5'd1, 4'd2, 4'd4, 16'd1942};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1942, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1720] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1721] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1722] = {5'd1, 4'd2, 4'd4, 16'd1943};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1943, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1723] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1724] = {5'd0, 4'd8, 4'd0, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 62, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1725] = {5'd1, 4'd2, 4'd4, 16'd1944};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1944, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1726] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1727] = {5'd0, 4'd8, 4'd0, 16'd108};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 108, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1728] = {5'd1, 4'd2, 4'd4, 16'd1945};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1945, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1729] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1730] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1731] = {5'd1, 4'd2, 4'd4, 16'd1946};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1946, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1732] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1733] = {5'd0, 4'd8, 4'd0, 16'd100};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 100, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1734] = {5'd1, 4'd2, 4'd4, 16'd1947};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1947, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1735] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1736] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1737] = {5'd1, 4'd2, 4'd4, 16'd1948};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1948, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1738] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1739] = {5'd0, 4'd8, 4'd0, 16'd52};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 52, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1740] = {5'd1, 4'd2, 4'd4, 16'd1949};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1949, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1741] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1742] = {5'd0, 4'd8, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 60, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1743] = {5'd1, 4'd2, 4'd4, 16'd1950};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1950, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1744] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1745] = {5'd0, 4'd8, 4'd0, 16'd47};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 47, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1746] = {5'd1, 4'd2, 4'd4, 16'd1951};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1951, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1747] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1748] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1749] = {5'd1, 4'd2, 4'd4, 16'd1952};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1952, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1750] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1751] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1752] = {5'd1, 4'd2, 4'd4, 16'd1953};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1953, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1753] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1754] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1755] = {5'd1, 4'd2, 4'd4, 16'd1954};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1954, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1756] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1757] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1758] = {5'd1, 4'd2, 4'd4, 16'd1955};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1955, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1759] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1760] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1761] = {5'd1, 4'd2, 4'd4, 16'd1956};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1956, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1762] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1763] = {5'd0, 4'd8, 4'd0, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 62, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1764] = {5'd1, 4'd2, 4'd4, 16'd1957};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1957, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1765] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1766] = {5'd0, 4'd8, 4'd0, 16'd9};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 9, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1767] = {5'd1, 4'd2, 4'd4, 16'd1958};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1958, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1768] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1769] = {5'd0, 4'd8, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 60, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1770] = {5'd1, 4'd2, 4'd4, 16'd1959};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1959, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1771] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1772] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1773] = {5'd1, 4'd2, 4'd4, 16'd1960};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1960, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1774] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1775] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1776] = {5'd1, 4'd2, 4'd4, 16'd1961};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1961, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1777] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1778] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1779] = {5'd1, 4'd2, 4'd4, 16'd1962};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1962, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1780] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1781] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1782] = {5'd1, 4'd2, 4'd4, 16'd1963};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1963, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1783] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1784] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1785] = {5'd1, 4'd2, 4'd4, 16'd1964};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1964, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1786] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1787] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1788] = {5'd1, 4'd2, 4'd4, 16'd1965};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1965, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1789] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1790] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1791] = {5'd1, 4'd2, 4'd4, 16'd1966};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1966, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1792] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1793] = {5'd0, 4'd8, 4'd0, 16'd121};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 121, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1794] = {5'd1, 4'd2, 4'd4, 16'd1967};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1967, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1795] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1796] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1797] = {5'd1, 4'd2, 4'd4, 16'd1968};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1968, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1798] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1799] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1800] = {5'd1, 4'd2, 4'd4, 16'd1969};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1969, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1801] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1802] = {5'd0, 4'd8, 4'd0, 16'd61};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 61, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1803] = {5'd1, 4'd2, 4'd4, 16'd1970};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1970, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1804] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1805] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1806] = {5'd1, 4'd2, 4'd4, 16'd1971};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1971, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1807] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1808] = {5'd0, 4'd8, 4'd0, 16'd99};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 99, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1809] = {5'd1, 4'd2, 4'd4, 16'd1972};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1972, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1810] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1811] = {5'd0, 4'd8, 4'd0, 16'd104};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 104, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1812] = {5'd1, 4'd2, 4'd4, 16'd1973};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1973, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1813] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1814] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1815] = {5'd1, 4'd2, 4'd4, 16'd1974};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1974, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1816] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1817] = {5'd0, 4'd8, 4'd0, 16'd99};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 99, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1818] = {5'd1, 4'd2, 4'd4, 16'd1975};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1975, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1819] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1820] = {5'd0, 4'd8, 4'd0, 16'd107};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 107, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1821] = {5'd1, 4'd2, 4'd4, 16'd1976};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1976, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1822] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1823] = {5'd0, 4'd8, 4'd0, 16'd98};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 98, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1824] = {5'd1, 4'd2, 4'd4, 16'd1977};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1977, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1825] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1826] = {5'd0, 4'd8, 4'd0, 16'd111};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 111, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1827] = {5'd1, 4'd2, 4'd4, 16'd1978};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1978, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1828] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1829] = {5'd0, 4'd8, 4'd0, 16'd120};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 120, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1830] = {5'd1, 4'd2, 4'd4, 16'd1979};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1979, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1831] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1832] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1833] = {5'd1, 4'd2, 4'd4, 16'd1980};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1980, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1834] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1835] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1836] = {5'd1, 4'd2, 4'd4, 16'd1981};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1981, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1837] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1838] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1839] = {5'd1, 4'd2, 4'd4, 16'd1982};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1982, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1840] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1841] = {5'd0, 4'd8, 4'd0, 16'd97};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 97, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1842] = {5'd1, 4'd2, 4'd4, 16'd1983};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1983, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1843] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1844] = {5'd0, 4'd8, 4'd0, 16'd109};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 109, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1845] = {5'd1, 4'd2, 4'd4, 16'd1984};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1984, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1846] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1847] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1848] = {5'd1, 4'd2, 4'd4, 16'd1985};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1985, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1849] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1850] = {5'd0, 4'd8, 4'd0, 16'd61};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 61, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1851] = {5'd1, 4'd2, 4'd4, 16'd1986};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1986, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1852] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1853] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1854] = {5'd1, 4'd2, 4'd4, 16'd1987};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1987, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1855] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1856] = {5'd0, 4'd8, 4'd0, 16'd108};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 108, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1857] = {5'd1, 4'd2, 4'd4, 16'd1988};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1988, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1858] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1859] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1860] = {5'd1, 4'd2, 4'd4, 16'd1989};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1989, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1861] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1862] = {5'd0, 4'd8, 4'd0, 16'd100};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 100, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1863] = {5'd1, 4'd2, 4'd4, 16'd1990};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1990, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1864] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1865] = {5'd0, 4'd8, 4'd0, 16'd52};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 52, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1866] = {5'd1, 4'd2, 4'd4, 16'd1991};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1991, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1867] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1868] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1869] = {5'd1, 4'd2, 4'd4, 16'd1992};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1992, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1870] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1871] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1872] = {5'd1, 4'd2, 4'd4, 16'd1993};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1993, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1873] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1874] = {5'd0, 4'd8, 4'd0, 16'd118};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 118, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1875] = {5'd1, 4'd2, 4'd4, 16'd1994};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1994, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1876] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1877] = {5'd0, 4'd8, 4'd0, 16'd97};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 97, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1878] = {5'd1, 4'd2, 4'd4, 16'd1995};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1995, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1879] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1880] = {5'd0, 4'd8, 4'd0, 16'd108};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 108, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1881] = {5'd1, 4'd2, 4'd4, 16'd1996};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1996, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1882] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1883] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1884] = {5'd1, 4'd2, 4'd4, 16'd1997};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1997, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1885] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1886] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1887] = {5'd1, 4'd2, 4'd4, 16'd1998};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1998, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1888] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1889] = {5'd0, 4'd8, 4'd0, 16'd61};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 61, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1890] = {5'd1, 4'd2, 4'd4, 16'd1999};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 1999, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1891] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1892] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1893] = {5'd1, 4'd2, 4'd4, 16'd2000};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2000, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1894] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1895] = {5'd0, 4'd8, 4'd0, 16'd70};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 70, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1896] = {5'd1, 4'd2, 4'd4, 16'd2001};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2001, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1897] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1898] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1899] = {5'd1, 4'd2, 4'd4, 16'd2002};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2002, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1900] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1901] = {5'd0, 4'd8, 4'd0, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 62, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1902] = {5'd1, 4'd2, 4'd4, 16'd2003};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2003, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1903] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1904] = {5'd0, 4'd8, 4'd0, 16'd108};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 108, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1905] = {5'd1, 4'd2, 4'd4, 16'd2004};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2004, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1906] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1907] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1908] = {5'd1, 4'd2, 4'd4, 16'd2005};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2005, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1909] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1910] = {5'd0, 4'd8, 4'd0, 16'd100};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 100, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1911] = {5'd1, 4'd2, 4'd4, 16'd2006};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2006, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1912] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1913] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1914] = {5'd1, 4'd2, 4'd4, 16'd2007};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2007, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1915] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1916] = {5'd0, 4'd8, 4'd0, 16'd53};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 53, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1917] = {5'd1, 4'd2, 4'd4, 16'd2008};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2008, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1918] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1919] = {5'd0, 4'd8, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 60, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1920] = {5'd1, 4'd2, 4'd4, 16'd2009};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2009, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1921] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1922] = {5'd0, 4'd8, 4'd0, 16'd47};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 47, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1923] = {5'd1, 4'd2, 4'd4, 16'd2010};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2010, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1924] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1925] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1926] = {5'd1, 4'd2, 4'd4, 16'd2011};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2011, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1927] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1928] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1929] = {5'd1, 4'd2, 4'd4, 16'd2012};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2012, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1930] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1931] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1932] = {5'd1, 4'd2, 4'd4, 16'd2013};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2013, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1933] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1934] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1935] = {5'd1, 4'd2, 4'd4, 16'd2014};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2014, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1936] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1937] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1938] = {5'd1, 4'd2, 4'd4, 16'd2015};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2015, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1939] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1940] = {5'd0, 4'd8, 4'd0, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 62, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1941] = {5'd1, 4'd2, 4'd4, 16'd2016};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2016, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1942] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1943] = {5'd0, 4'd8, 4'd0, 16'd9};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 9, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1944] = {5'd1, 4'd2, 4'd4, 16'd2017};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2017, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1945] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1946] = {5'd0, 4'd8, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 60, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1947] = {5'd1, 4'd2, 4'd4, 16'd2018};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2018, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1948] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1949] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1950] = {5'd1, 4'd2, 4'd4, 16'd2019};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2019, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1951] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1952] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1953] = {5'd1, 4'd2, 4'd4, 16'd2020};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2020, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1954] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1955] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1956] = {5'd1, 4'd2, 4'd4, 16'd2021};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2021, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1957] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1958] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1959] = {5'd1, 4'd2, 4'd4, 16'd2022};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2022, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1960] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1961] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1962] = {5'd1, 4'd2, 4'd4, 16'd2023};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2023, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1963] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1964] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1965] = {5'd1, 4'd2, 4'd4, 16'd2024};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2024, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1966] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1967] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1968] = {5'd1, 4'd2, 4'd4, 16'd2025};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2025, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1969] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1970] = {5'd0, 4'd8, 4'd0, 16'd121};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 121, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1971] = {5'd1, 4'd2, 4'd4, 16'd2026};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2026, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1972] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1973] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1974] = {5'd1, 4'd2, 4'd4, 16'd2027};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2027, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1975] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1976] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1977] = {5'd1, 4'd2, 4'd4, 16'd2028};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2028, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1978] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1979] = {5'd0, 4'd8, 4'd0, 16'd61};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 61, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1980] = {5'd1, 4'd2, 4'd4, 16'd2029};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2029, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1981] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1982] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1983] = {5'd1, 4'd2, 4'd4, 16'd2030};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2030, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1984] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1985] = {5'd0, 4'd8, 4'd0, 16'd99};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 99, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1986] = {5'd1, 4'd2, 4'd4, 16'd2031};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2031, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1987] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1988] = {5'd0, 4'd8, 4'd0, 16'd104};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 104, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1989] = {5'd1, 4'd2, 4'd4, 16'd2032};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2032, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1990] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1991] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1992] = {5'd1, 4'd2, 4'd4, 16'd2033};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2033, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1993] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1994] = {5'd0, 4'd8, 4'd0, 16'd99};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 99, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1995] = {5'd1, 4'd2, 4'd4, 16'd2034};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2034, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1996] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[1997] = {5'd0, 4'd8, 4'd0, 16'd107};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 107, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[1998] = {5'd1, 4'd2, 4'd4, 16'd2035};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2035, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[1999] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2000] = {5'd0, 4'd8, 4'd0, 16'd98};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 98, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2001] = {5'd1, 4'd2, 4'd4, 16'd2036};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2036, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2002] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2003] = {5'd0, 4'd8, 4'd0, 16'd111};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 111, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2004] = {5'd1, 4'd2, 4'd4, 16'd2037};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2037, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2005] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2006] = {5'd0, 4'd8, 4'd0, 16'd120};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 120, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2007] = {5'd1, 4'd2, 4'd4, 16'd2038};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2038, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2008] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2009] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2010] = {5'd1, 4'd2, 4'd4, 16'd2039};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2039, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2011] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2012] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2013] = {5'd1, 4'd2, 4'd4, 16'd2040};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2040, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2014] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2015] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2016] = {5'd1, 4'd2, 4'd4, 16'd2041};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2041, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2017] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2018] = {5'd0, 4'd8, 4'd0, 16'd97};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 97, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2019] = {5'd1, 4'd2, 4'd4, 16'd2042};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2042, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2020] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2021] = {5'd0, 4'd8, 4'd0, 16'd109};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 109, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2022] = {5'd1, 4'd2, 4'd4, 16'd2043};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2043, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2023] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2024] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2025] = {5'd1, 4'd2, 4'd4, 16'd2044};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2044, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2026] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2027] = {5'd0, 4'd8, 4'd0, 16'd61};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 61, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2028] = {5'd1, 4'd2, 4'd4, 16'd2045};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2045, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2029] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2030] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2031] = {5'd1, 4'd2, 4'd4, 16'd2046};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2046, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2032] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2033] = {5'd0, 4'd8, 4'd0, 16'd108};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 108, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2034] = {5'd1, 4'd2, 4'd4, 16'd2047};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2047, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2035] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2036] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2037] = {5'd1, 4'd2, 4'd4, 16'd2048};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2048, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2038] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2039] = {5'd0, 4'd8, 4'd0, 16'd100};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 100, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2040] = {5'd1, 4'd2, 4'd4, 16'd2049};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2049, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2041] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2042] = {5'd0, 4'd8, 4'd0, 16'd52};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 52, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2043] = {5'd1, 4'd2, 4'd4, 16'd2050};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2050, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2044] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2045] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2046] = {5'd1, 4'd2, 4'd4, 16'd2051};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2051, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2047] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2048] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2049] = {5'd1, 4'd2, 4'd4, 16'd2052};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2052, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2050] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2051] = {5'd0, 4'd8, 4'd0, 16'd118};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 118, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2052] = {5'd1, 4'd2, 4'd4, 16'd2053};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2053, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2053] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2054] = {5'd0, 4'd8, 4'd0, 16'd97};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 97, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2055] = {5'd1, 4'd2, 4'd4, 16'd2054};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2054, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2056] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2057] = {5'd0, 4'd8, 4'd0, 16'd108};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 108, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2058] = {5'd1, 4'd2, 4'd4, 16'd2055};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2055, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2059] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2060] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2061] = {5'd1, 4'd2, 4'd4, 16'd2056};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2056, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2062] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2063] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2064] = {5'd1, 4'd2, 4'd4, 16'd2057};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2057, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2065] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2066] = {5'd0, 4'd8, 4'd0, 16'd61};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 61, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2067] = {5'd1, 4'd2, 4'd4, 16'd2058};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2058, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2068] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2069] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2070] = {5'd1, 4'd2, 4'd4, 16'd2059};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2059, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2071] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2072] = {5'd0, 4'd8, 4'd0, 16'd71};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 71, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2073] = {5'd1, 4'd2, 4'd4, 16'd2060};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2060, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2074] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2075] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2076] = {5'd1, 4'd2, 4'd4, 16'd2061};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2061, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2077] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2078] = {5'd0, 4'd8, 4'd0, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 62, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2079] = {5'd1, 4'd2, 4'd4, 16'd2062};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2062, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2080] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2081] = {5'd0, 4'd8, 4'd0, 16'd108};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 108, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2082] = {5'd1, 4'd2, 4'd4, 16'd2063};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2063, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2083] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2084] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2085] = {5'd1, 4'd2, 4'd4, 16'd2064};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2064, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2086] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2087] = {5'd0, 4'd8, 4'd0, 16'd100};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 100, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2088] = {5'd1, 4'd2, 4'd4, 16'd2065};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2065, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2089] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2090] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2091] = {5'd1, 4'd2, 4'd4, 16'd2066};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2066, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2092] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2093] = {5'd0, 4'd8, 4'd0, 16'd54};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 54, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2094] = {5'd1, 4'd2, 4'd4, 16'd2067};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2067, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2095] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2096] = {5'd0, 4'd8, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 60, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2097] = {5'd1, 4'd2, 4'd4, 16'd2068};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2068, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2098] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2099] = {5'd0, 4'd8, 4'd0, 16'd47};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 47, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2100] = {5'd1, 4'd2, 4'd4, 16'd2069};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2069, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2101] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2102] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2103] = {5'd1, 4'd2, 4'd4, 16'd2070};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2070, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2104] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2105] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2106] = {5'd1, 4'd2, 4'd4, 16'd2071};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2071, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2107] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2108] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2109] = {5'd1, 4'd2, 4'd4, 16'd2072};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2072, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2110] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2111] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2112] = {5'd1, 4'd2, 4'd4, 16'd2073};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2073, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2113] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2114] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2115] = {5'd1, 4'd2, 4'd4, 16'd2074};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2074, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2116] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2117] = {5'd0, 4'd8, 4'd0, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 62, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2118] = {5'd1, 4'd2, 4'd4, 16'd2075};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2075, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2119] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2120] = {5'd0, 4'd8, 4'd0, 16'd9};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 9, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2121] = {5'd1, 4'd2, 4'd4, 16'd2076};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2076, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2122] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2123] = {5'd0, 4'd8, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 60, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2124] = {5'd1, 4'd2, 4'd4, 16'd2077};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2077, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2125] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2126] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2127] = {5'd1, 4'd2, 4'd4, 16'd2078};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2078, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2128] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2129] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2130] = {5'd1, 4'd2, 4'd4, 16'd2079};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2079, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2131] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2132] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2133] = {5'd1, 4'd2, 4'd4, 16'd2080};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2080, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2134] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2135] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2136] = {5'd1, 4'd2, 4'd4, 16'd2081};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2081, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2137] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2138] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2139] = {5'd1, 4'd2, 4'd4, 16'd2082};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2082, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2140] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2141] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2142] = {5'd1, 4'd2, 4'd4, 16'd2083};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2083, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2143] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2144] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2145] = {5'd1, 4'd2, 4'd4, 16'd2084};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2084, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2146] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2147] = {5'd0, 4'd8, 4'd0, 16'd121};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 121, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2148] = {5'd1, 4'd2, 4'd4, 16'd2085};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2085, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2149] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2150] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2151] = {5'd1, 4'd2, 4'd4, 16'd2086};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2086, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2152] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2153] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2154] = {5'd1, 4'd2, 4'd4, 16'd2087};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2087, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2155] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2156] = {5'd0, 4'd8, 4'd0, 16'd61};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 61, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2157] = {5'd1, 4'd2, 4'd4, 16'd2088};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2088, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2158] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2159] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2160] = {5'd1, 4'd2, 4'd4, 16'd2089};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2089, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2161] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2162] = {5'd0, 4'd8, 4'd0, 16'd99};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 99, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2163] = {5'd1, 4'd2, 4'd4, 16'd2090};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2090, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2164] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2165] = {5'd0, 4'd8, 4'd0, 16'd104};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 104, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2166] = {5'd1, 4'd2, 4'd4, 16'd2091};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2091, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2167] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2168] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2169] = {5'd1, 4'd2, 4'd4, 16'd2092};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2092, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2170] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2171] = {5'd0, 4'd8, 4'd0, 16'd99};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 99, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2172] = {5'd1, 4'd2, 4'd4, 16'd2093};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2093, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2173] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2174] = {5'd0, 4'd8, 4'd0, 16'd107};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 107, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2175] = {5'd1, 4'd2, 4'd4, 16'd2094};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2094, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2176] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2177] = {5'd0, 4'd8, 4'd0, 16'd98};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 98, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2178] = {5'd1, 4'd2, 4'd4, 16'd2095};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2095, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2179] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2180] = {5'd0, 4'd8, 4'd0, 16'd111};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 111, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2181] = {5'd1, 4'd2, 4'd4, 16'd2096};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2096, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2182] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2183] = {5'd0, 4'd8, 4'd0, 16'd120};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 120, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2184] = {5'd1, 4'd2, 4'd4, 16'd2097};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2097, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2185] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2186] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2187] = {5'd1, 4'd2, 4'd4, 16'd2098};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2098, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2188] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2189] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2190] = {5'd1, 4'd2, 4'd4, 16'd2099};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2099, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2191] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2192] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2193] = {5'd1, 4'd2, 4'd4, 16'd2100};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2100, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2194] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2195] = {5'd0, 4'd8, 4'd0, 16'd97};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 97, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2196] = {5'd1, 4'd2, 4'd4, 16'd2101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2101, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2197] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2198] = {5'd0, 4'd8, 4'd0, 16'd109};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 109, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2199] = {5'd1, 4'd2, 4'd4, 16'd2102};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2102, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2200] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2201] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2202] = {5'd1, 4'd2, 4'd4, 16'd2103};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2103, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2203] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2204] = {5'd0, 4'd8, 4'd0, 16'd61};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 61, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2205] = {5'd1, 4'd2, 4'd4, 16'd2104};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2104, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2206] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2207] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2208] = {5'd1, 4'd2, 4'd4, 16'd2105};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2105, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2209] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2210] = {5'd0, 4'd8, 4'd0, 16'd108};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 108, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2211] = {5'd1, 4'd2, 4'd4, 16'd2106};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2106, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2212] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2213] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2214] = {5'd1, 4'd2, 4'd4, 16'd2107};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2107, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2215] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2216] = {5'd0, 4'd8, 4'd0, 16'd100};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 100, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2217] = {5'd1, 4'd2, 4'd4, 16'd2108};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2108, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2218] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2219] = {5'd0, 4'd8, 4'd0, 16'd52};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 52, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2220] = {5'd1, 4'd2, 4'd4, 16'd2109};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2109, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2221] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2222] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2223] = {5'd1, 4'd2, 4'd4, 16'd2110};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2110, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2224] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2225] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2226] = {5'd1, 4'd2, 4'd4, 16'd2111};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2111, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2227] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2228] = {5'd0, 4'd8, 4'd0, 16'd118};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 118, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2229] = {5'd1, 4'd2, 4'd4, 16'd2112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2112, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2230] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2231] = {5'd0, 4'd8, 4'd0, 16'd97};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 97, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2232] = {5'd1, 4'd2, 4'd4, 16'd2113};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2113, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2233] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2234] = {5'd0, 4'd8, 4'd0, 16'd108};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 108, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2235] = {5'd1, 4'd2, 4'd4, 16'd2114};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2114, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2236] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2237] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2238] = {5'd1, 4'd2, 4'd4, 16'd2115};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2115, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2239] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2240] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2241] = {5'd1, 4'd2, 4'd4, 16'd2116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2116, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2242] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2243] = {5'd0, 4'd8, 4'd0, 16'd61};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 61, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2244] = {5'd1, 4'd2, 4'd4, 16'd2117};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2117, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2245] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2246] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2247] = {5'd1, 4'd2, 4'd4, 16'd2118};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2118, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2248] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2249] = {5'd0, 4'd8, 4'd0, 16'd72};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 72, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2250] = {5'd1, 4'd2, 4'd4, 16'd2119};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2119, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2251] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2252] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2253] = {5'd1, 4'd2, 4'd4, 16'd2120};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2120, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2254] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2255] = {5'd0, 4'd8, 4'd0, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 62, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2256] = {5'd1, 4'd2, 4'd4, 16'd2121};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2121, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2257] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2258] = {5'd0, 4'd8, 4'd0, 16'd108};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 108, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2259] = {5'd1, 4'd2, 4'd4, 16'd2122};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2122, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2260] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2261] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2262] = {5'd1, 4'd2, 4'd4, 16'd2123};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2123, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2263] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2264] = {5'd0, 4'd8, 4'd0, 16'd100};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 100, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2265] = {5'd1, 4'd2, 4'd4, 16'd2124};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2124, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2266] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2267] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2268] = {5'd1, 4'd2, 4'd4, 16'd2125};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2125, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2269] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2270] = {5'd0, 4'd8, 4'd0, 16'd55};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 55, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2271] = {5'd1, 4'd2, 4'd4, 16'd2126};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2126, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2272] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2273] = {5'd0, 4'd8, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 60, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2274] = {5'd1, 4'd2, 4'd4, 16'd2127};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2127, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2275] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2276] = {5'd0, 4'd8, 4'd0, 16'd47};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 47, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2277] = {5'd1, 4'd2, 4'd4, 16'd2128};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2128, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2278] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2279] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2280] = {5'd1, 4'd2, 4'd4, 16'd2129};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2129, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2281] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2282] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2283] = {5'd1, 4'd2, 4'd4, 16'd2130};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2130, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2284] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2285] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2286] = {5'd1, 4'd2, 4'd4, 16'd2131};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2131, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2287] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2288] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2289] = {5'd1, 4'd2, 4'd4, 16'd2132};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2132, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2290] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2291] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2292] = {5'd1, 4'd2, 4'd4, 16'd2133};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2133, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2293] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2294] = {5'd0, 4'd8, 4'd0, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 62, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2295] = {5'd1, 4'd2, 4'd4, 16'd2134};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2134, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2296] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2297] = {5'd0, 4'd8, 4'd0, 16'd9};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 9, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2298] = {5'd1, 4'd2, 4'd4, 16'd2135};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2135, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2299] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2300] = {5'd0, 4'd8, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 60, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2301] = {5'd1, 4'd2, 4'd4, 16'd2136};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2136, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2302] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2303] = {5'd0, 4'd8, 4'd0, 16'd98};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 98, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2304] = {5'd1, 4'd2, 4'd4, 16'd2137};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2137, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2305] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2306] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2307] = {5'd1, 4'd2, 4'd4, 16'd2138};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2138, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2308] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2309] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2310] = {5'd1, 4'd2, 4'd4, 16'd2139};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2139, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2311] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2312] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2313] = {5'd1, 4'd2, 4'd4, 16'd2140};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2140, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2314] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2315] = {5'd0, 4'd8, 4'd0, 16'd111};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 111, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2316] = {5'd1, 4'd2, 4'd4, 16'd2141};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2141, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2317] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2318] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2319] = {5'd1, 4'd2, 4'd4, 16'd2142};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2142, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2320] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2321] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2322] = {5'd1, 4'd2, 4'd4, 16'd2143};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2143, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2323] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2324] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2325] = {5'd1, 4'd2, 4'd4, 16'd2144};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2144, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2326] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2327] = {5'd0, 4'd8, 4'd0, 16'd121};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 121, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2328] = {5'd1, 4'd2, 4'd4, 16'd2145};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2145, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2329] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2330] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2331] = {5'd1, 4'd2, 4'd4, 16'd2146};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2146, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2332] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2333] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2334] = {5'd1, 4'd2, 4'd4, 16'd2147};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2147, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2335] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2336] = {5'd0, 4'd8, 4'd0, 16'd61};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 61, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2337] = {5'd1, 4'd2, 4'd4, 16'd2148};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2148, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2338] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2339] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2340] = {5'd1, 4'd2, 4'd4, 16'd2149};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2149, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2341] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2342] = {5'd0, 4'd8, 4'd0, 16'd115};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 115, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2343] = {5'd1, 4'd2, 4'd4, 16'd2150};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2150, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2344] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2345] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2346] = {5'd1, 4'd2, 4'd4, 16'd2151};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2151, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2347] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2348] = {5'd0, 4'd8, 4'd0, 16'd109};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 109, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2349] = {5'd1, 4'd2, 4'd4, 16'd2152};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2152, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2350] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2351] = {5'd0, 4'd8, 4'd0, 16'd98};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 98, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2352] = {5'd1, 4'd2, 4'd4, 16'd2153};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2153, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2353] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2354] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2355] = {5'd1, 4'd2, 4'd4, 16'd2154};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2154, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2356] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2357] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2358] = {5'd1, 4'd2, 4'd4, 16'd2155};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2155, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2359] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2360] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2361] = {5'd1, 4'd2, 4'd4, 16'd2156};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2156, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2362] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2363] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2364] = {5'd1, 4'd2, 4'd4, 16'd2157};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2157, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2365] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2366] = {5'd0, 4'd8, 4'd0, 16'd118};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 118, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2367] = {5'd1, 4'd2, 4'd4, 16'd2158};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2158, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2368] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2369] = {5'd0, 4'd8, 4'd0, 16'd97};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 97, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2370] = {5'd1, 4'd2, 4'd4, 16'd2159};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2159, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2371] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2372] = {5'd0, 4'd8, 4'd0, 16'd108};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 108, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2373] = {5'd1, 4'd2, 4'd4, 16'd2160};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2160, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2374] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2375] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2376] = {5'd1, 4'd2, 4'd4, 16'd2161};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2161, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2377] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2378] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2379] = {5'd1, 4'd2, 4'd4, 16'd2162};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2162, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2380] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2381] = {5'd0, 4'd8, 4'd0, 16'd61};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 61, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2382] = {5'd1, 4'd2, 4'd4, 16'd2163};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2163, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2383] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2384] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2385] = {5'd1, 4'd2, 4'd4, 16'd2164};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2164, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2386] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2387] = {5'd0, 4'd8, 4'd0, 16'd83};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 83, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2388] = {5'd1, 4'd2, 4'd4, 16'd2165};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2165, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2389] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2390] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2391] = {5'd1, 4'd2, 4'd4, 16'd2166};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2166, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2392] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2393] = {5'd0, 4'd8, 4'd0, 16'd98};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 98, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2394] = {5'd1, 4'd2, 4'd4, 16'd2167};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2167, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2395] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2396] = {5'd0, 4'd8, 4'd0, 16'd109};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 109, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2397] = {5'd1, 4'd2, 4'd4, 16'd2168};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2168, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2398] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2399] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2400] = {5'd1, 4'd2, 4'd4, 16'd2169};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2169, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2401] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2402] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2403] = {5'd1, 4'd2, 4'd4, 16'd2170};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2170, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2404] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2405] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2406] = {5'd1, 4'd2, 4'd4, 16'd2171};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2171, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2407] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2408] = {5'd0, 4'd8, 4'd0, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 62, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2409] = {5'd1, 4'd2, 4'd4, 16'd2172};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2172, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2410] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2411] = {5'd0, 4'd8, 4'd0, 16'd85};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 85, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2412] = {5'd1, 4'd2, 4'd4, 16'd2173};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2173, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2413] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2414] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2415] = {5'd1, 4'd2, 4'd4, 16'd2174};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2174, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2416] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2417] = {5'd0, 4'd8, 4'd0, 16'd100};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 100, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2418] = {5'd1, 4'd2, 4'd4, 16'd2175};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2175, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2419] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2420] = {5'd0, 4'd8, 4'd0, 16'd97};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 97, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2421] = {5'd1, 4'd2, 4'd4, 16'd2176};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2176, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2422] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2423] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2424] = {5'd1, 4'd2, 4'd4, 16'd2177};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2177, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2425] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2426] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2427] = {5'd1, 4'd2, 4'd4, 16'd2178};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2178, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2428] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2429] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2430] = {5'd1, 4'd2, 4'd4, 16'd2179};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2179, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2431] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2432] = {5'd0, 4'd8, 4'd0, 16'd76};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 76, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2433] = {5'd1, 4'd2, 4'd4, 16'd2180};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2180, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2434] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2435] = {5'd0, 4'd8, 4'd0, 16'd69};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 69, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2436] = {5'd1, 4'd2, 4'd4, 16'd2181};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2181, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2437] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2438] = {5'd0, 4'd8, 4'd0, 16'd68};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 68, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2439] = {5'd1, 4'd2, 4'd4, 16'd2182};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2182, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2440] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2441] = {5'd0, 4'd8, 4'd0, 16'd115};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 115, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2442] = {5'd1, 4'd2, 4'd4, 16'd2183};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2183, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2443] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2444] = {5'd0, 4'd8, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 60, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2445] = {5'd1, 4'd2, 4'd4, 16'd2184};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2184, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2446] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2447] = {5'd0, 4'd8, 4'd0, 16'd47};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 47, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2448] = {5'd1, 4'd2, 4'd4, 16'd2185};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2185, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2449] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2450] = {5'd0, 4'd8, 4'd0, 16'd98};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 98, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2451] = {5'd1, 4'd2, 4'd4, 16'd2186};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2186, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2452] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2453] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2454] = {5'd1, 4'd2, 4'd4, 16'd2187};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2187, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2455] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2456] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2457] = {5'd1, 4'd2, 4'd4, 16'd2188};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2188, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2458] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2459] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2460] = {5'd1, 4'd2, 4'd4, 16'd2189};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2189, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2461] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2462] = {5'd0, 4'd8, 4'd0, 16'd111};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 111, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2463] = {5'd1, 4'd2, 4'd4, 16'd2190};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2190, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2464] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2465] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2466] = {5'd1, 4'd2, 4'd4, 16'd2191};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2191, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2467] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2468] = {5'd0, 4'd8, 4'd0, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 62, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2469] = {5'd1, 4'd2, 4'd4, 16'd2192};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2192, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2470] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2471] = {5'd0, 4'd8, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 60, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2472] = {5'd1, 4'd2, 4'd4, 16'd2193};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2193, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2473] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2474] = {5'd0, 4'd8, 4'd0, 16'd47};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 47, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2475] = {5'd1, 4'd2, 4'd4, 16'd2194};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2194, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2476] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2477] = {5'd0, 4'd8, 4'd0, 16'd102};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 102, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2478] = {5'd1, 4'd2, 4'd4, 16'd2195};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2195, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2479] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2480] = {5'd0, 4'd8, 4'd0, 16'd111};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 111, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2481] = {5'd1, 4'd2, 4'd4, 16'd2196};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2196, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2482] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2483] = {5'd0, 4'd8, 4'd0, 16'd114};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 114, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2484] = {5'd1, 4'd2, 4'd4, 16'd2197};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2197, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2485] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2486] = {5'd0, 4'd8, 4'd0, 16'd109};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 109, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2487] = {5'd1, 4'd2, 4'd4, 16'd2198};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2198, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2488] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2489] = {5'd0, 4'd8, 4'd0, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 62, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2490] = {5'd1, 4'd2, 4'd4, 16'd2199};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2199, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2491] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2492] = {5'd0, 4'd8, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 60, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2493] = {5'd1, 4'd2, 4'd4, 16'd2200};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2200, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2494] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2495] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2496] = {5'd1, 4'd2, 4'd4, 16'd2201};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2201, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2497] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2498] = {5'd0, 4'd8, 4'd0, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 62, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2499] = {5'd1, 4'd2, 4'd4, 16'd2202};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2202, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2500] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2501] = {5'd0, 4'd8, 4'd0, 16'd84};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 84, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2502] = {5'd1, 4'd2, 4'd4, 16'd2203};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2203, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2503] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2504] = {5'd0, 4'd8, 4'd0, 16'd104};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 104, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2505] = {5'd1, 4'd2, 4'd4, 16'd2204};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2204, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2506] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2507] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2508] = {5'd1, 4'd2, 4'd4, 16'd2205};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2205, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2509] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2510] = {5'd0, 4'd8, 4'd0, 16'd115};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 115, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2511] = {5'd1, 4'd2, 4'd4, 16'd2206};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2206, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2512] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2513] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2514] = {5'd1, 4'd2, 4'd4, 16'd2207};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2207, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2515] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2516] = {5'd0, 4'd8, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 60, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2517] = {5'd1, 4'd2, 4'd4, 16'd2208};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2208, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2518] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2519] = {5'd0, 4'd8, 4'd0, 16'd97};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 97, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2520] = {5'd1, 4'd2, 4'd4, 16'd2209};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2209, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2521] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2522] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2523] = {5'd1, 4'd2, 4'd4, 16'd2210};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2210, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2524] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2525] = {5'd0, 4'd8, 4'd0, 16'd104};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 104, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2526] = {5'd1, 4'd2, 4'd4, 16'd2211};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2211, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2527] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2528] = {5'd0, 4'd8, 4'd0, 16'd114};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 114, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2529] = {5'd1, 4'd2, 4'd4, 16'd2212};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2212, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2530] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2531] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2532] = {5'd1, 4'd2, 4'd4, 16'd2213};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2213, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2533] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2534] = {5'd0, 4'd8, 4'd0, 16'd102};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 102, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2535] = {5'd1, 4'd2, 4'd4, 16'd2214};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2214, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2536] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2537] = {5'd0, 4'd8, 4'd0, 16'd61};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 61, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2538] = {5'd1, 4'd2, 4'd4, 16'd2215};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2215, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2539] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2540] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2541] = {5'd1, 4'd2, 4'd4, 16'd2216};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2216, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2542] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2543] = {5'd0, 4'd8, 4'd0, 16'd104};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 104, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2544] = {5'd1, 4'd2, 4'd4, 16'd2217};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2217, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2545] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2546] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2547] = {5'd1, 4'd2, 4'd4, 16'd2218};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2218, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2548] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2549] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2550] = {5'd1, 4'd2, 4'd4, 16'd2219};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2219, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2551] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2552] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2553] = {5'd1, 4'd2, 4'd4, 16'd2220};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2220, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2554] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2555] = {5'd0, 4'd8, 4'd0, 16'd115};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 115, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2556] = {5'd1, 4'd2, 4'd4, 16'd2221};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2221, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2557] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2558] = {5'd0, 4'd8, 4'd0, 16'd58};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 58, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2559] = {5'd1, 4'd2, 4'd4, 16'd2222};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2222, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2560] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2561] = {5'd0, 4'd8, 4'd0, 16'd47};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 47, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2562] = {5'd1, 4'd2, 4'd4, 16'd2223};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2223, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2563] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2564] = {5'd0, 4'd8, 4'd0, 16'd47};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 47, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2565] = {5'd1, 4'd2, 4'd4, 16'd2224};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2224, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2566] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2567] = {5'd0, 4'd8, 4'd0, 16'd103};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 103, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2568] = {5'd1, 4'd2, 4'd4, 16'd2225};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2225, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2569] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2570] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2571] = {5'd1, 4'd2, 4'd4, 16'd2226};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2226, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2572] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2573] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2574] = {5'd1, 4'd2, 4'd4, 16'd2227};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2227, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2575] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2576] = {5'd0, 4'd8, 4'd0, 16'd104};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 104, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2577] = {5'd1, 4'd2, 4'd4, 16'd2228};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2228, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2578] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2579] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2580] = {5'd1, 4'd2, 4'd4, 16'd2229};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2229, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2581] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2582] = {5'd0, 4'd8, 4'd0, 16'd98};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 98, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2583] = {5'd1, 4'd2, 4'd4, 16'd2230};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2230, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2584] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2585] = {5'd0, 4'd8, 4'd0, 16'd46};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 46, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2586] = {5'd1, 4'd2, 4'd4, 16'd2231};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2231, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2587] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2588] = {5'd0, 4'd8, 4'd0, 16'd99};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 99, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2589] = {5'd1, 4'd2, 4'd4, 16'd2232};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2232, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2590] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2591] = {5'd0, 4'd8, 4'd0, 16'd111};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 111, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2592] = {5'd1, 4'd2, 4'd4, 16'd2233};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2233, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2593] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2594] = {5'd0, 4'd8, 4'd0, 16'd109};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 109, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2595] = {5'd1, 4'd2, 4'd4, 16'd2234};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2234, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2596] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2597] = {5'd0, 4'd8, 4'd0, 16'd47};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 47, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2598] = {5'd1, 4'd2, 4'd4, 16'd2235};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2235, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2599] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2600] = {5'd0, 4'd8, 4'd0, 16'd100};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 100, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2601] = {5'd1, 4'd2, 4'd4, 16'd2236};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2236, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2602] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2603] = {5'd0, 4'd8, 4'd0, 16'd97};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 97, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2604] = {5'd1, 4'd2, 4'd4, 16'd2237};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2237, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2605] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2606] = {5'd0, 4'd8, 4'd0, 16'd119};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 119, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2607] = {5'd1, 4'd2, 4'd4, 16'd2238};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2238, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2608] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2609] = {5'd0, 4'd8, 4'd0, 16'd115};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 115, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2610] = {5'd1, 4'd2, 4'd4, 16'd2239};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2239, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2611] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2612] = {5'd0, 4'd8, 4'd0, 16'd111};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 111, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2613] = {5'd1, 4'd2, 4'd4, 16'd2240};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2240, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2614] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2615] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2616] = {5'd1, 4'd2, 4'd4, 16'd2241};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2241, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2617] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2618] = {5'd0, 4'd8, 4'd0, 16'd106};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 106, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2619] = {5'd1, 4'd2, 4'd4, 16'd2242};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2242, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2620] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2621] = {5'd0, 4'd8, 4'd0, 16'd111};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 111, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2622] = {5'd1, 4'd2, 4'd4, 16'd2243};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2243, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2623] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2624] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2625] = {5'd1, 4'd2, 4'd4, 16'd2244};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2244, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2626] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2627] = {5'd0, 4'd8, 4'd0, 16'd47};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 47, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2628] = {5'd1, 4'd2, 4'd4, 16'd2245};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2245, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2629] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2630] = {5'd0, 4'd8, 4'd0, 16'd67};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 67, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2631] = {5'd1, 4'd2, 4'd4, 16'd2246};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2246, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2632] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2633] = {5'd0, 4'd8, 4'd0, 16'd104};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 104, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2634] = {5'd1, 4'd2, 4'd4, 16'd2247};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2247, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2635] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2636] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2637] = {5'd1, 4'd2, 4'd4, 16'd2248};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2248, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2638] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2639] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2640] = {5'd1, 4'd2, 4'd4, 16'd2249};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2249, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2641] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2642] = {5'd0, 4'd8, 4'd0, 16'd115};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 115, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2643] = {5'd1, 4'd2, 4'd4, 16'd2250};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2250, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2644] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2645] = {5'd0, 4'd8, 4'd0, 16'd45};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 45, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2646] = {5'd1, 4'd2, 4'd4, 16'd2251};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2251, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2647] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2648] = {5'd0, 4'd8, 4'd0, 16'd68};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 68, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2649] = {5'd1, 4'd2, 4'd4, 16'd2252};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2252, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2650] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2651] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2652] = {5'd1, 4'd2, 4'd4, 16'd2253};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2253, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2653] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2654] = {5'd0, 4'd8, 4'd0, 16'd109};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 109, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2655] = {5'd1, 4'd2, 4'd4, 16'd2254};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2254, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2656] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2657] = {5'd0, 4'd8, 4'd0, 16'd111};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 111, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2658] = {5'd1, 4'd2, 4'd4, 16'd2255};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2255, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2659] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2660] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2661] = {5'd1, 4'd2, 4'd4, 16'd2256};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2256, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2662] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2663] = {5'd0, 4'd8, 4'd0, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 62, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2664] = {5'd1, 4'd2, 4'd4, 16'd2257};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2257, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2665] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2666] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2667] = {5'd1, 4'd2, 4'd4, 16'd2258};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2258, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2668] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2669] = {5'd0, 4'd8, 4'd0, 16'd114};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 114, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2670] = {5'd1, 4'd2, 4'd4, 16'd2259};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2259, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2671] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2672] = {5'd0, 4'd8, 4'd0, 16'd111};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 111, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2673] = {5'd1, 4'd2, 4'd4, 16'd2260};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2260, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2674] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2675] = {5'd0, 4'd8, 4'd0, 16'd106};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 106, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2676] = {5'd1, 4'd2, 4'd4, 16'd2261};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2261, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2677] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2678] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2679] = {5'd1, 4'd2, 4'd4, 16'd2262};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2262, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2680] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2681] = {5'd0, 4'd8, 4'd0, 16'd99};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 99, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2682] = {5'd1, 4'd2, 4'd4, 16'd2263};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2263, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2683] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2684] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2685] = {5'd1, 4'd2, 4'd4, 16'd2264};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2264, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2686] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2687] = {5'd0, 4'd8, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 60, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2688] = {5'd1, 4'd2, 4'd4, 16'd2265};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2265, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2689] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2690] = {5'd0, 4'd8, 4'd0, 16'd47};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 47, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2691] = {5'd1, 4'd2, 4'd4, 16'd2266};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2266, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2692] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2693] = {5'd0, 4'd8, 4'd0, 16'd97};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 97, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2694] = {5'd1, 4'd2, 4'd4, 16'd2267};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2267, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2695] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2696] = {5'd0, 4'd8, 4'd0, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 62, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2697] = {5'd1, 4'd2, 4'd4, 16'd2268};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2268, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2698] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2699] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2700] = {5'd1, 4'd2, 4'd4, 16'd2269};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2269, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2701] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2702] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2703] = {5'd1, 4'd2, 4'd4, 16'd2270};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2270, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2704] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2705] = {5'd0, 4'd8, 4'd0, 16'd115};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 115, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2706] = {5'd1, 4'd2, 4'd4, 16'd2271};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2271, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2707] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2708] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2709] = {5'd1, 4'd2, 4'd4, 16'd2272};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2272, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2710] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2711] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2712] = {5'd1, 4'd2, 4'd4, 16'd2273};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2273, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2713] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2714] = {5'd0, 4'd8, 4'd0, 16'd111};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 111, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2715] = {5'd1, 4'd2, 4'd4, 16'd2274};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2274, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2716] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2717] = {5'd0, 4'd8, 4'd0, 16'd119};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 119, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2718] = {5'd1, 4'd2, 4'd4, 16'd2275};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2275, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2719] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2720] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2721] = {5'd1, 4'd2, 4'd4, 16'd2276};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2276, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2722] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2723] = {5'd0, 4'd8, 4'd0, 16'd114};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 114, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2724] = {5'd1, 4'd2, 4'd4, 16'd2277};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2277, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2725] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2726] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2727] = {5'd1, 4'd2, 4'd4, 16'd2278};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2278, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2728] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2729] = {5'd0, 4'd8, 4'd0, 16'd100};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 100, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2730] = {5'd1, 4'd2, 4'd4, 16'd2279};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2279, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2731] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2732] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2733] = {5'd1, 4'd2, 4'd4, 16'd2280};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2280, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2734] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2735] = {5'd0, 4'd8, 4'd0, 16'd98};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 98, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2736] = {5'd1, 4'd2, 4'd4, 16'd2281};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2281, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2737] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2738] = {5'd0, 4'd8, 4'd0, 16'd121};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 121, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2739] = {5'd1, 4'd2, 4'd4, 16'd2282};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2282, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2740] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2741] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2742] = {5'd1, 4'd2, 4'd4, 16'd2283};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2283, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2743] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2744] = {5'd0, 4'd8, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 60, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2745] = {5'd1, 4'd2, 4'd4, 16'd2284};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2284, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2746] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2747] = {5'd0, 4'd8, 4'd0, 16'd97};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 97, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2748] = {5'd1, 4'd2, 4'd4, 16'd2285};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2285, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2749] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2750] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2751] = {5'd1, 4'd2, 4'd4, 16'd2286};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2286, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2752] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2753] = {5'd0, 4'd8, 4'd0, 16'd104};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 104, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2754] = {5'd1, 4'd2, 4'd4, 16'd2287};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2287, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2755] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2756] = {5'd0, 4'd8, 4'd0, 16'd114};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 114, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2757] = {5'd1, 4'd2, 4'd4, 16'd2288};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2288, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2758] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2759] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2760] = {5'd1, 4'd2, 4'd4, 16'd2289};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2289, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2761] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2762] = {5'd0, 4'd8, 4'd0, 16'd102};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 102, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2763] = {5'd1, 4'd2, 4'd4, 16'd2290};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2290, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2764] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2765] = {5'd0, 4'd8, 4'd0, 16'd61};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 61, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2766] = {5'd1, 4'd2, 4'd4, 16'd2291};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2291, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2767] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2768] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2769] = {5'd1, 4'd2, 4'd4, 16'd2292};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2292, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2770] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2771] = {5'd0, 4'd8, 4'd0, 16'd104};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 104, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2772] = {5'd1, 4'd2, 4'd4, 16'd2293};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2293, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2773] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2774] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2775] = {5'd1, 4'd2, 4'd4, 16'd2294};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2294, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2776] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2777] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2778] = {5'd1, 4'd2, 4'd4, 16'd2295};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2295, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2779] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2780] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2781] = {5'd1, 4'd2, 4'd4, 16'd2296};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2296, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2782] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2783] = {5'd0, 4'd8, 4'd0, 16'd58};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 58, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2784] = {5'd1, 4'd2, 4'd4, 16'd2297};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2297, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2785] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2786] = {5'd0, 4'd8, 4'd0, 16'd47};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 47, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2787] = {5'd1, 4'd2, 4'd4, 16'd2298};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2298, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2788] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2789] = {5'd0, 4'd8, 4'd0, 16'd47};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 47, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2790] = {5'd1, 4'd2, 4'd4, 16'd2299};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2299, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2791] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2792] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2793] = {5'd1, 4'd2, 4'd4, 16'd2300};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2300, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2794] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2795] = {5'd0, 4'd8, 4'd0, 16'd121};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 121, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2796] = {5'd1, 4'd2, 4'd4, 16'd2301};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2301, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2797] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2798] = {5'd0, 4'd8, 4'd0, 16'd97};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 97, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2799] = {5'd1, 4'd2, 4'd4, 16'd2302};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2302, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2800] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2801] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2802] = {5'd1, 4'd2, 4'd4, 16'd2303};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2303, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2803] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2804] = {5'd0, 4'd8, 4'd0, 16'd100};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 100, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2805] = {5'd1, 4'd2, 4'd4, 16'd2304};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2304, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2806] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2807] = {5'd0, 4'd8, 4'd0, 16'd99};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 99, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2808] = {5'd1, 4'd2, 4'd4, 16'd2305};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2305, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2809] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2810] = {5'd0, 4'd8, 4'd0, 16'd104};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 104, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2811] = {5'd1, 4'd2, 4'd4, 16'd2306};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2306, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2812] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2813] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2814] = {5'd1, 4'd2, 4'd4, 16'd2307};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2307, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2815] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2816] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2817] = {5'd1, 4'd2, 4'd4, 16'd2308};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2308, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2818] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2819] = {5'd0, 4'd8, 4'd0, 16'd115};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 115, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2820] = {5'd1, 4'd2, 4'd4, 16'd2309};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2309, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2821] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2822] = {5'd0, 4'd8, 4'd0, 16'd46};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 46, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2823] = {5'd1, 4'd2, 4'd4, 16'd2310};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2310, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2824] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2825] = {5'd0, 4'd8, 4'd0, 16'd111};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 111, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2826] = {5'd1, 4'd2, 4'd4, 16'd2311};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2311, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2827] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2828] = {5'd0, 4'd8, 4'd0, 16'd114};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 114, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2829] = {5'd1, 4'd2, 4'd4, 16'd2312};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2312, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2830] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2831] = {5'd0, 4'd8, 4'd0, 16'd103};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 103, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2832] = {5'd1, 4'd2, 4'd4, 16'd2313};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2313, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2833] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2834] = {5'd0, 4'd8, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 34, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2835] = {5'd1, 4'd2, 4'd4, 16'd2314};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2314, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2836] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2837] = {5'd0, 4'd8, 4'd0, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 62, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2838] = {5'd1, 4'd2, 4'd4, 16'd2315};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2315, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2839] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2840] = {5'd0, 4'd8, 4'd0, 16'd67};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 67, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2841] = {5'd1, 4'd2, 4'd4, 16'd2316};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2316, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2842] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2843] = {5'd0, 4'd8, 4'd0, 16'd104};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 104, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2844] = {5'd1, 4'd2, 4'd4, 16'd2317};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2317, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2845] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2846] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2847] = {5'd1, 4'd2, 4'd4, 16'd2318};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2318, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2848] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2849] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2850] = {5'd1, 4'd2, 4'd4, 16'd2319};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2319, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2851] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2852] = {5'd0, 4'd8, 4'd0, 16'd115};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 115, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2853] = {5'd1, 4'd2, 4'd4, 16'd2320};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2320, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2854] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2855] = {5'd0, 4'd8, 4'd0, 16'd45};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 45, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2856] = {5'd1, 4'd2, 4'd4, 16'd2321};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2321, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2857] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2858] = {5'd0, 4'd8, 4'd0, 16'd50};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 50, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2859] = {5'd1, 4'd2, 4'd4, 16'd2322};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2322, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2860] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2861] = {5'd0, 4'd8, 4'd0, 16'd46};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 46, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2862] = {5'd1, 4'd2, 4'd4, 16'd2323};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2323, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2863] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2864] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2865] = {5'd1, 4'd2, 4'd4, 16'd2324};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2324, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2866] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2867] = {5'd0, 4'd8, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 60, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2868] = {5'd1, 4'd2, 4'd4, 16'd2325};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2325, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2869] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2870] = {5'd0, 4'd8, 4'd0, 16'd47};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 47, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2871] = {5'd1, 4'd2, 4'd4, 16'd2326};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2326, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2872] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2873] = {5'd0, 4'd8, 4'd0, 16'd97};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 97, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2874] = {5'd1, 4'd2, 4'd4, 16'd2327};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2327, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2875] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2876] = {5'd0, 4'd8, 4'd0, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 62, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2877] = {5'd1, 4'd2, 4'd4, 16'd2328};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2328, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2878] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2879] = {5'd0, 4'd8, 4'd0, 16'd46};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 46, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2880] = {5'd1, 4'd2, 4'd4, 16'd2329};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2329, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2881] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2882] = {5'd0, 4'd8, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 60, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2883] = {5'd1, 4'd2, 4'd4, 16'd2330};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2330, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2884] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2885] = {5'd0, 4'd8, 4'd0, 16'd47};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 47, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2886] = {5'd1, 4'd2, 4'd4, 16'd2331};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2331, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2887] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2888] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2889] = {5'd1, 4'd2, 4'd4, 16'd2332};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2332, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2890] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2891] = {5'd0, 4'd8, 4'd0, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 62, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2892] = {5'd1, 4'd2, 4'd4, 16'd2333};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2333, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2893] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2894] = {5'd0, 4'd8, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 60, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2895] = {5'd1, 4'd2, 4'd4, 16'd2334};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2334, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2896] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2897] = {5'd0, 4'd8, 4'd0, 16'd47};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 47, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2898] = {5'd1, 4'd2, 4'd4, 16'd2335};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2335, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2899] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2900] = {5'd0, 4'd8, 4'd0, 16'd98};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 98, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2901] = {5'd1, 4'd2, 4'd4, 16'd2336};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2336, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2902] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2903] = {5'd0, 4'd8, 4'd0, 16'd111};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 111, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2904] = {5'd1, 4'd2, 4'd4, 16'd2337};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2337, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2905] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2906] = {5'd0, 4'd8, 4'd0, 16'd100};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 100, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2907] = {5'd1, 4'd2, 4'd4, 16'd2338};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2338, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2908] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2909] = {5'd0, 4'd8, 4'd0, 16'd121};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 121, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2910] = {5'd1, 4'd2, 4'd4, 16'd2339};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2339, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2911] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2912] = {5'd0, 4'd8, 4'd0, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 62, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2913] = {5'd1, 4'd2, 4'd4, 16'd2340};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2340, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2914] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2915] = {5'd0, 4'd8, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 60, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2916] = {5'd1, 4'd2, 4'd4, 16'd2341};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2341, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2917] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2918] = {5'd0, 4'd8, 4'd0, 16'd47};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 47, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2919] = {5'd1, 4'd2, 4'd4, 16'd2342};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2342, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2920] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2921] = {5'd0, 4'd8, 4'd0, 16'd104};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 104, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2922] = {5'd1, 4'd2, 4'd4, 16'd2343};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2343, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2923] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2924] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2925] = {5'd1, 4'd2, 4'd4, 16'd2344};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2344, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2926] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2927] = {5'd0, 4'd8, 4'd0, 16'd109};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 109, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2928] = {5'd1, 4'd2, 4'd4, 16'd2345};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2345, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2929] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2930] = {5'd0, 4'd8, 4'd0, 16'd108};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 108, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2931] = {5'd1, 4'd2, 4'd4, 16'd2346};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2346, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2932] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2933] = {5'd0, 4'd8, 4'd0, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 62, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2934] = {5'd1, 4'd2, 4'd4, 16'd2347};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2347, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2935] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2936] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'literal'}
    instructions[2937] = {5'd1, 4'd2, 4'd4, 16'd2348};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 4, 'literal': 2348, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'addl'}
    instructions[2938] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 62, 'op': 'store'}
    instructions[2939] = {5'd0, 4'd8, 4'd0, 16'd52};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 87 {'literal': 52, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 87, 'op': 'literal'}
    instructions[2940] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 87 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 87, 'op': 'addl'}
    instructions[2941] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 87 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 87, 'op': 'load'}
    instructions[2942] = {5'd0, 4'd2, 4'd0, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 87 {'literal': 7, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 87, 'op': 'literal'}
    instructions[2943] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 87 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 87, 'op': 'store'}
    instructions[2944] = {5'd0, 4'd8, 4'd0, 16'd50};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 88 {'literal': 50, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 88, 'op': 'literal'}
    instructions[2945] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 88 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 88, 'op': 'addl'}
    instructions[2946] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 88 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 88, 'op': 'load'}
    instructions[2947] = {5'd0, 4'd2, 4'd0, 16'd9};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 88 {'literal': 9, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 88, 'op': 'literal'}
    instructions[2948] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 88 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 88, 'op': 'store'}
    instructions[2949] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'store'}
    instructions[2950] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'addl'}
    instructions[2951] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'store'}
    instructions[2952] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'addl'}
    instructions[2953] = {5'd0, 4'd8, 4'd0, 16'd12};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'literal': 12, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'literal'}
    instructions[2954] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'store'}
    instructions[2955] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'addl'}
    instructions[2956] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'addl'}
    instructions[2957] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'addl'}
    instructions[2958] = {5'd3, 4'd6, 4'd0, 16'd4497};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'z': 6, 'label': 4497, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'call'}
    instructions[2959] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'addl'}
    instructions[2960] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2961] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'load'}
    instructions[2962] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2963] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'load'}
    instructions[2964] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 90, 'op': 'addl'}
    instructions[2965] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'store'}
    instructions[2966] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'addl'}
    instructions[2967] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'store'}
    instructions[2968] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'addl'}
    instructions[2969] = {5'd0, 4'd8, 4'd0, 16'd54};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'literal': 54, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'literal'}
    instructions[2970] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'store'}
    instructions[2971] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'addl'}
    instructions[2972] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'addl'}
    instructions[2973] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'addl'}
    instructions[2974] = {5'd3, 4'd6, 4'd0, 16'd4497};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'z': 6, 'label': 4497, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'call'}
    instructions[2975] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'addl'}
    instructions[2976] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2977] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'load'}
    instructions[2978] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2979] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'load'}
    instructions[2980] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 91, 'op': 'addl'}
    instructions[2981] = {5'd0, 4'd8, 4'd0, 16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 94 {'literal': 5, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 94, 'op': 'literal'}
    instructions[2982] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 94 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 94, 'op': 'addl'}
    instructions[2983] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 94 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 94, 'op': 'load'}
    instructions[2984] = {5'd6, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 94 {'a': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 94, 'op': 'read'}
    instructions[2985] = {5'd1, 4'd2, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 94 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 94, 'op': 'addl'}
    instructions[2986] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 94 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 94, 'op': 'store'}
    instructions[2987] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 95 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 95, 'op': 'literal'}
    instructions[2988] = {5'd1, 4'd2, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 95 {'a': 4, 'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 95, 'op': 'addl'}
    instructions[2989] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 95 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 95, 'op': 'store'}
    instructions[2990] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96, 'op': 'literal'}
    instructions[2991] = {5'd1, 4'd2, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96 {'a': 4, 'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96, 'op': 'addl'}
    instructions[2992] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96, 'op': 'store'}
    instructions[2993] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96, 'op': 'addl'}
    instructions[2994] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96, 'op': 'addl'}
    instructions[2995] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96, 'op': 'load'}
    instructions[2996] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96, 'op': 'store'}
    instructions[2997] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96, 'op': 'addl'}
    instructions[2998] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96, 'op': 'addl'}
    instructions[2999] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96, 'op': 'addl'}
    instructions[3000] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96, 'op': 'load'}
    instructions[3001] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3002] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96, 'op': 'load'}
    instructions[3003] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96, 'op': 'unsigned_greater'}
    instructions[3004] = {5'd8, 4'd0, 4'd8, 16'd3113};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96 {'a': 8, 'label': 3113, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96, 'op': 'jmp_if_false'}
    instructions[3005] = {5'd0, 4'd8, 4'd0, 16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 97 {'literal': 5, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 97, 'op': 'literal'}
    instructions[3006] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 97 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 97, 'op': 'addl'}
    instructions[3007] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 97 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 97, 'op': 'load'}
    instructions[3008] = {5'd6, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 97 {'a': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 97, 'op': 'read'}
    instructions[3009] = {5'd1, 4'd2, 4'd4, 16'd1463};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 97 {'a': 4, 'literal': 1463, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 97, 'op': 'addl'}
    instructions[3010] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 97 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 97, 'op': 'store'}
    instructions[3011] = {5'd0, 4'd8, 4'd0, 16'd255};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98 {'literal': 255, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98, 'op': 'literal'}
    instructions[3012] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98, 'op': 'store'}
    instructions[3013] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98, 'op': 'addl'}
    instructions[3014] = {5'd0, 4'd8, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98 {'literal': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98, 'op': 'literal'}
    instructions[3015] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98, 'op': 'store'}
    instructions[3016] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98, 'op': 'addl'}
    instructions[3017] = {5'd1, 4'd8, 4'd4, 16'd1463};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98 {'a': 4, 'literal': 1463, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98, 'op': 'addl'}
    instructions[3018] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98, 'op': 'addl'}
    instructions[3019] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98, 'op': 'load'}
    instructions[3020] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3021] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98, 'op': 'load'}
    instructions[3022] = {5'd9, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98, 'op': 'unsigned_shift_right'}
    instructions[3023] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3024] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98, 'op': 'load'}
    instructions[3025] = {5'd10, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98, 'op': 'and'}
    instructions[3026] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98, 'op': 'store'}
    instructions[3027] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98, 'op': 'addl'}
    instructions[3028] = {5'd1, 4'd8, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98 {'a': 4, 'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98, 'op': 'addl'}
    instructions[3029] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98, 'op': 'store'}
    instructions[3030] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98, 'op': 'addl'}
    instructions[3031] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98, 'op': 'addl'}
    instructions[3032] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98, 'op': 'addl'}
    instructions[3033] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98, 'op': 'load'}
    instructions[3034] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3035] = {5'd5, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98, 'op': 'load'}
    instructions[3036] = {5'd11, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98, 'op': 'add'}
    instructions[3037] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98, 'op': 'addl'}
    instructions[3038] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3039] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98, 'op': 'load'}
    instructions[3040] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 98, 'op': 'store'}
    instructions[3041] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 99 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 99, 'op': 'addl'}
    instructions[3042] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 99 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 99, 'op': 'addl'}
    instructions[3043] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 99 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 99, 'op': 'load'}
    instructions[3044] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 99 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 99, 'op': 'store'}
    instructions[3045] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 99 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 99, 'op': 'addl'}
    instructions[3046] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 99 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 99, 'op': 'literal'}
    instructions[3047] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 99 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 99, 'op': 'store'}
    instructions[3048] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 99 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 99, 'op': 'addl'}
    instructions[3049] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 99 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 99, 'op': 'addl'}
    instructions[3050] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 99 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 99, 'op': 'addl'}
    instructions[3051] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 99 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 99, 'op': 'load'}
    instructions[3052] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 99 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 99, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3053] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 99 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 99, 'op': 'load'}
    instructions[3054] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 99 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 99, 'op': 'add'}
    instructions[3055] = {5'd1, 4'd2, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 99 {'a': 4, 'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 99, 'op': 'addl'}
    instructions[3056] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 99 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 99, 'op': 'store'}
    instructions[3057] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 99 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 99, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3058] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 99 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 99, 'op': 'load'}
    instructions[3059] = {5'd0, 4'd8, 4'd0, 16'd255};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100 {'literal': 255, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100, 'op': 'literal'}
    instructions[3060] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100, 'op': 'store'}
    instructions[3061] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100, 'op': 'addl'}
    instructions[3062] = {5'd1, 4'd8, 4'd4, 16'd1463};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100 {'a': 4, 'literal': 1463, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100, 'op': 'addl'}
    instructions[3063] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100, 'op': 'addl'}
    instructions[3064] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100, 'op': 'load'}
    instructions[3065] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3066] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100, 'op': 'load'}
    instructions[3067] = {5'd10, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100, 'op': 'and'}
    instructions[3068] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100, 'op': 'store'}
    instructions[3069] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100, 'op': 'addl'}
    instructions[3070] = {5'd1, 4'd8, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100 {'a': 4, 'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100, 'op': 'addl'}
    instructions[3071] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100, 'op': 'store'}
    instructions[3072] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100, 'op': 'addl'}
    instructions[3073] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100, 'op': 'addl'}
    instructions[3074] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100, 'op': 'addl'}
    instructions[3075] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100, 'op': 'load'}
    instructions[3076] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3077] = {5'd5, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100, 'op': 'load'}
    instructions[3078] = {5'd11, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100, 'op': 'add'}
    instructions[3079] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100, 'op': 'addl'}
    instructions[3080] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3081] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100, 'op': 'load'}
    instructions[3082] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 100, 'op': 'store'}
    instructions[3083] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 101 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 101, 'op': 'addl'}
    instructions[3084] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 101 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 101, 'op': 'addl'}
    instructions[3085] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 101 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 101, 'op': 'load'}
    instructions[3086] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 101 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 101, 'op': 'store'}
    instructions[3087] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 101 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 101, 'op': 'addl'}
    instructions[3088] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 101 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 101, 'op': 'literal'}
    instructions[3089] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 101 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 101, 'op': 'store'}
    instructions[3090] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 101 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 101, 'op': 'addl'}
    instructions[3091] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 101 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 101, 'op': 'addl'}
    instructions[3092] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 101 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 101, 'op': 'addl'}
    instructions[3093] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 101 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 101, 'op': 'load'}
    instructions[3094] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 101 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 101, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3095] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 101 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 101, 'op': 'load'}
    instructions[3096] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 101 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 101, 'op': 'add'}
    instructions[3097] = {5'd1, 4'd2, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 101 {'a': 4, 'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 101, 'op': 'addl'}
    instructions[3098] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 101 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 101, 'op': 'store'}
    instructions[3099] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 101 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 101, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3100] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 101 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 101, 'op': 'load'}
    instructions[3101] = {5'd0, 4'd8, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96 {'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96, 'op': 'literal'}
    instructions[3102] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96, 'op': 'store'}
    instructions[3103] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96, 'op': 'addl'}
    instructions[3104] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96, 'op': 'addl'}
    instructions[3105] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96, 'op': 'addl'}
    instructions[3106] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96, 'op': 'load'}
    instructions[3107] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3108] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96, 'op': 'load'}
    instructions[3109] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96, 'op': 'add'}
    instructions[3110] = {5'd1, 4'd2, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96 {'a': 4, 'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96, 'op': 'addl'}
    instructions[3111] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96, 'op': 'store'}
    instructions[3112] = {5'd12, 4'd0, 4'd0, 16'd2993};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96 {'label': 2993, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 96, 'op': 'goto'}
    instructions[3113] = {5'd0, 4'd8, 4'd0, 16'd71};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 107 {'literal': 71, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 107, 'op': 'literal'}
    instructions[3114] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 107 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 107, 'op': 'store'}
    instructions[3115] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 107 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 107, 'op': 'addl'}
    instructions[3116] = {5'd1, 4'd8, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 107 {'a': 4, 'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 107, 'op': 'addl'}
    instructions[3117] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 107 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 107, 'op': 'store'}
    instructions[3118] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 107 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 107, 'op': 'addl'}
    instructions[3119] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 107 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 107, 'op': 'literal'}
    instructions[3120] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 107 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 107, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3121] = {5'd5, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 107 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 107, 'op': 'load'}
    instructions[3122] = {5'd11, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 107 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 107, 'op': 'add'}
    instructions[3123] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 107 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 107, 'op': 'addl'}
    instructions[3124] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 107 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 107, 'op': 'load'}
    instructions[3125] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 107 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 107, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3126] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 107 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 107, 'op': 'load'}
    instructions[3127] = {5'd13, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 107 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 107, 'op': 'equal'}
    instructions[3128] = {5'd8, 4'd0, 4'd8, 16'd3144};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 108 {'a': 8, 'label': 3144, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 108, 'op': 'jmp_if_false'}
    instructions[3129] = {5'd0, 4'd8, 4'd0, 16'd69};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 108 {'literal': 69, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 108, 'op': 'literal'}
    instructions[3130] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 108 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 108, 'op': 'store'}
    instructions[3131] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 108 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 108, 'op': 'addl'}
    instructions[3132] = {5'd1, 4'd8, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 108 {'a': 4, 'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 108, 'op': 'addl'}
    instructions[3133] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 108 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 108, 'op': 'store'}
    instructions[3134] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 108 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 108, 'op': 'addl'}
    instructions[3135] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 108 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 108, 'op': 'literal'}
    instructions[3136] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 108 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 108, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3137] = {5'd5, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 108 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 108, 'op': 'load'}
    instructions[3138] = {5'd11, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 108 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 108, 'op': 'add'}
    instructions[3139] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 108 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 108, 'op': 'addl'}
    instructions[3140] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 108 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 108, 'op': 'load'}
    instructions[3141] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 108 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 108, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3142] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 108 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 108, 'op': 'load'}
    instructions[3143] = {5'd13, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 108 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 108, 'op': 'equal'}
    instructions[3144] = {5'd8, 4'd0, 4'd8, 16'd3160};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 109 {'a': 8, 'label': 3160, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 109, 'op': 'jmp_if_false'}
    instructions[3145] = {5'd0, 4'd8, 4'd0, 16'd84};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 109 {'literal': 84, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 109, 'op': 'literal'}
    instructions[3146] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 109 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 109, 'op': 'store'}
    instructions[3147] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 109 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 109, 'op': 'addl'}
    instructions[3148] = {5'd1, 4'd8, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 109 {'a': 4, 'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 109, 'op': 'addl'}
    instructions[3149] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 109 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 109, 'op': 'store'}
    instructions[3150] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 109 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 109, 'op': 'addl'}
    instructions[3151] = {5'd0, 4'd8, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 109 {'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 109, 'op': 'literal'}
    instructions[3152] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 109 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 109, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3153] = {5'd5, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 109 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 109, 'op': 'load'}
    instructions[3154] = {5'd11, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 109 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 109, 'op': 'add'}
    instructions[3155] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 109 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 109, 'op': 'addl'}
    instructions[3156] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 109 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 109, 'op': 'load'}
    instructions[3157] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 109 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 109, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3158] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 109 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 109, 'op': 'load'}
    instructions[3159] = {5'd13, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 109 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 109, 'op': 'equal'}
    instructions[3160] = {5'd8, 4'd0, 4'd8, 16'd3176};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 110 {'a': 8, 'label': 3176, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 110, 'op': 'jmp_if_false'}
    instructions[3161] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 110 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 110, 'op': 'literal'}
    instructions[3162] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 110 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 110, 'op': 'store'}
    instructions[3163] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 110 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 110, 'op': 'addl'}
    instructions[3164] = {5'd1, 4'd8, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 110 {'a': 4, 'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 110, 'op': 'addl'}
    instructions[3165] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 110 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 110, 'op': 'store'}
    instructions[3166] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 110 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 110, 'op': 'addl'}
    instructions[3167] = {5'd0, 4'd8, 4'd0, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 110 {'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 110, 'op': 'literal'}
    instructions[3168] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 110 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 110, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3169] = {5'd5, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 110 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 110, 'op': 'load'}
    instructions[3170] = {5'd11, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 110 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 110, 'op': 'add'}
    instructions[3171] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 110 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 110, 'op': 'addl'}
    instructions[3172] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 110 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 110, 'op': 'load'}
    instructions[3173] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 110 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 110, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3174] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 110 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 110, 'op': 'load'}
    instructions[3175] = {5'd13, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 110 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 110, 'op': 'equal'}
    instructions[3176] = {5'd8, 4'd0, 4'd8, 16'd3192};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 111 {'a': 8, 'label': 3192, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 111, 'op': 'jmp_if_false'}
    instructions[3177] = {5'd0, 4'd8, 4'd0, 16'd47};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 111 {'literal': 47, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 111, 'op': 'literal'}
    instructions[3178] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 111 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 111, 'op': 'store'}
    instructions[3179] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 111 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 111, 'op': 'addl'}
    instructions[3180] = {5'd1, 4'd8, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 111 {'a': 4, 'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 111, 'op': 'addl'}
    instructions[3181] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 111 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 111, 'op': 'store'}
    instructions[3182] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 111 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 111, 'op': 'addl'}
    instructions[3183] = {5'd0, 4'd8, 4'd0, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 111 {'literal': 4, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 111, 'op': 'literal'}
    instructions[3184] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 111 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 111, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3185] = {5'd5, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 111 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 111, 'op': 'load'}
    instructions[3186] = {5'd11, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 111 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 111, 'op': 'add'}
    instructions[3187] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 111 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 111, 'op': 'addl'}
    instructions[3188] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 111 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 111, 'op': 'load'}
    instructions[3189] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 111 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 111, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3190] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 111 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 111, 'op': 'load'}
    instructions[3191] = {5'd13, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 111 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 111, 'op': 'equal'}
    instructions[3192] = {5'd8, 4'd0, 4'd8, 16'd3224};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112 {'a': 8, 'label': 3224, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112, 'op': 'jmp_if_false'}
    instructions[3193] = {5'd0, 4'd8, 4'd0, 16'd63};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112 {'literal': 63, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112, 'op': 'literal'}
    instructions[3194] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112, 'op': 'store'}
    instructions[3195] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112, 'op': 'addl'}
    instructions[3196] = {5'd1, 4'd8, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112 {'a': 4, 'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112, 'op': 'addl'}
    instructions[3197] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112, 'op': 'store'}
    instructions[3198] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112, 'op': 'addl'}
    instructions[3199] = {5'd0, 4'd8, 4'd0, 16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112 {'literal': 5, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112, 'op': 'literal'}
    instructions[3200] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3201] = {5'd5, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112, 'op': 'load'}
    instructions[3202] = {5'd11, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112, 'op': 'add'}
    instructions[3203] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112, 'op': 'addl'}
    instructions[3204] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112, 'op': 'load'}
    instructions[3205] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3206] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112, 'op': 'load'}
    instructions[3207] = {5'd13, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112, 'op': 'equal'}
    instructions[3208] = {5'd14, 4'd0, 4'd8, 16'd3224};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112 {'a': 8, 'label': 3224, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112, 'op': 'jmp_if_true'}
    instructions[3209] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112, 'op': 'literal'}
    instructions[3210] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112, 'op': 'store'}
    instructions[3211] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112, 'op': 'addl'}
    instructions[3212] = {5'd1, 4'd8, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112 {'a': 4, 'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112, 'op': 'addl'}
    instructions[3213] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112, 'op': 'store'}
    instructions[3214] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112, 'op': 'addl'}
    instructions[3215] = {5'd0, 4'd8, 4'd0, 16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112 {'literal': 5, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112, 'op': 'literal'}
    instructions[3216] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3217] = {5'd5, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112, 'op': 'load'}
    instructions[3218] = {5'd11, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112, 'op': 'add'}
    instructions[3219] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112, 'op': 'addl'}
    instructions[3220] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112, 'op': 'load'}
    instructions[3221] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3222] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112, 'op': 'load'}
    instructions[3223] = {5'd13, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 112, 'op': 'equal'}
    instructions[3224] = {5'd8, 4'd0, 4'd8, 16'd4480};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 107 {'a': 8, 'label': 4480, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 107, 'op': 'jmp_if_false'}
    instructions[3225] = {5'd0, 4'd8, 4'd0, 16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 113 {'literal': 5, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 113, 'op': 'literal'}
    instructions[3226] = {5'd1, 4'd2, 4'd4, 16'd1467};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 113 {'a': 4, 'literal': 1467, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 113, 'op': 'addl'}
    instructions[3227] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 113 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 113, 'op': 'store'}
    instructions[3228] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114, 'op': 'store'}
    instructions[3229] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114, 'op': 'addl'}
    instructions[3230] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114, 'op': 'store'}
    instructions[3231] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114, 'op': 'addl'}
    instructions[3232] = {5'd1, 4'd8, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114 {'a': 4, 'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114, 'op': 'addl'}
    instructions[3233] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114, 'op': 'store'}
    instructions[3234] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114, 'op': 'addl'}
    instructions[3235] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114, 'op': 'literal'}
    instructions[3236] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114, 'op': 'store'}
    instructions[3237] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114, 'op': 'addl'}
    instructions[3238] = {5'd1, 4'd8, 4'd4, 16'd1467};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114 {'a': 4, 'literal': 1467, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114, 'op': 'addl'}
    instructions[3239] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114, 'op': 'addl'}
    instructions[3240] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114, 'op': 'load'}
    instructions[3241] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114, 'op': 'store'}
    instructions[3242] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114, 'op': 'addl'}
    instructions[3243] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114, 'op': 'addl'}
    instructions[3244] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114, 'op': 'addl'}
    instructions[3245] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114, 'op': 'load'}
    instructions[3246] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114, 'op': 'store'}
    instructions[3247] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114, 'op': 'addl'}
    instructions[3248] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114, 'op': 'addl'}
    instructions[3249] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114, 'op': 'addl'}
    instructions[3250] = {5'd3, 4'd6, 4'd0, 16'd4588};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114 {'z': 6, 'label': 4588, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114, 'op': 'call'}
    instructions[3251] = {5'd1, 4'd3, 4'd3, -16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114 {'a': 3, 'literal': -4, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114, 'op': 'addl'}
    instructions[3252] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3253] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114, 'op': 'load'}
    instructions[3254] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3255] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114, 'op': 'load'}
    instructions[3256] = {5'd0, 4'd2, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114 {'literal': 6, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114, 'op': 'literal'}
    instructions[3257] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114, 'op': 'load'}
    instructions[3258] = {5'd1, 4'd2, 4'd4, 16'd1468};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114 {'a': 4, 'literal': 1468, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114, 'op': 'addl'}
    instructions[3259] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 114, 'op': 'store'}
    instructions[3260] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 115 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 115, 'op': 'literal'}
    instructions[3261] = {5'd1, 4'd2, 4'd4, 16'd1466};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 115 {'a': 4, 'literal': 1466, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 115, 'op': 'addl'}
    instructions[3262] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 115 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 115, 'op': 'store'}
    instructions[3263] = {5'd0, 4'd8, 4'd0, 16'd65535};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'literal': 65535, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'op': 'literal'}
    instructions[3264] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'op': 'store'}
    instructions[3265] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'op': 'addl'}
    instructions[3266] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'op': 'store'}
    instructions[3267] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'op': 'addl'}
    instructions[3268] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'op': 'store'}
    instructions[3269] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'op': 'addl'}
    instructions[3270] = {5'd1, 4'd8, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'a': 4, 'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'op': 'addl'}
    instructions[3271] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'op': 'store'}
    instructions[3272] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'op': 'addl'}
    instructions[3273] = {5'd0, 4'd8, 4'd0, 16'd65};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'literal': 65, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'op': 'literal'}
    instructions[3274] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'op': 'store'}
    instructions[3275] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'op': 'addl'}
    instructions[3276] = {5'd1, 4'd8, 4'd4, 16'd1467};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'a': 4, 'literal': 1467, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'op': 'addl'}
    instructions[3277] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'op': 'addl'}
    instructions[3278] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'op': 'load'}
    instructions[3279] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'op': 'store'}
    instructions[3280] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'op': 'addl'}
    instructions[3281] = {5'd1, 4'd8, 4'd4, 16'd1468};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'a': 4, 'literal': 1468, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'op': 'addl'}
    instructions[3282] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'op': 'addl'}
    instructions[3283] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'op': 'load'}
    instructions[3284] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'op': 'store'}
    instructions[3285] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'op': 'addl'}
    instructions[3286] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'op': 'addl'}
    instructions[3287] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'op': 'addl'}
    instructions[3288] = {5'd3, 4'd6, 4'd0, 16'd4588};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'z': 6, 'label': 4588, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'op': 'call'}
    instructions[3289] = {5'd1, 4'd3, 4'd3, -16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'a': 3, 'literal': -4, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'op': 'addl'}
    instructions[3290] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3291] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'op': 'load'}
    instructions[3292] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3293] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'op': 'load'}
    instructions[3294] = {5'd0, 4'd2, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'literal': 6, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'op': 'literal'}
    instructions[3295] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'op': 'load'}
    instructions[3296] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3297] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'op': 'load'}
    instructions[3298] = {5'd15, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'op': 'not_equal'}
    instructions[3299] = {5'd8, 4'd0, 4'd8, 16'd3312};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'a': 8, 'label': 3312, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'op': 'jmp_if_false'}
    instructions[3300] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'op': 'literal'}
    instructions[3301] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'op': 'store'}
    instructions[3302] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'op': 'addl'}
    instructions[3303] = {5'd1, 4'd8, 4'd4, 16'd1466};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'a': 4, 'literal': 1466, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'op': 'addl'}
    instructions[3304] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'op': 'addl'}
    instructions[3305] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'op': 'load'}
    instructions[3306] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3307] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'op': 'load'}
    instructions[3308] = {5'd16, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'op': 'or'}
    instructions[3309] = {5'd1, 4'd2, 4'd4, 16'd1466};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'a': 4, 'literal': 1466, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'op': 'addl'}
    instructions[3310] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'op': 'store'}
    instructions[3311] = {5'd12, 4'd0, 4'd0, 16'd3312};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116 {'label': 3312, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 116, 'op': 'goto'}
    instructions[3312] = {5'd0, 4'd8, 4'd0, 16'd65535};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'literal': 65535, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'op': 'literal'}
    instructions[3313] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'op': 'store'}
    instructions[3314] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'op': 'addl'}
    instructions[3315] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'op': 'store'}
    instructions[3316] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'op': 'addl'}
    instructions[3317] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'op': 'store'}
    instructions[3318] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'op': 'addl'}
    instructions[3319] = {5'd1, 4'd8, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'a': 4, 'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'op': 'addl'}
    instructions[3320] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'op': 'store'}
    instructions[3321] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'op': 'addl'}
    instructions[3322] = {5'd0, 4'd8, 4'd0, 16'd66};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'literal': 66, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'op': 'literal'}
    instructions[3323] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'op': 'store'}
    instructions[3324] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'op': 'addl'}
    instructions[3325] = {5'd1, 4'd8, 4'd4, 16'd1467};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'a': 4, 'literal': 1467, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'op': 'addl'}
    instructions[3326] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'op': 'addl'}
    instructions[3327] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'op': 'load'}
    instructions[3328] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'op': 'store'}
    instructions[3329] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'op': 'addl'}
    instructions[3330] = {5'd1, 4'd8, 4'd4, 16'd1468};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'a': 4, 'literal': 1468, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'op': 'addl'}
    instructions[3331] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'op': 'addl'}
    instructions[3332] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'op': 'load'}
    instructions[3333] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'op': 'store'}
    instructions[3334] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'op': 'addl'}
    instructions[3335] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'op': 'addl'}
    instructions[3336] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'op': 'addl'}
    instructions[3337] = {5'd3, 4'd6, 4'd0, 16'd4588};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'z': 6, 'label': 4588, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'op': 'call'}
    instructions[3338] = {5'd1, 4'd3, 4'd3, -16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'a': 3, 'literal': -4, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'op': 'addl'}
    instructions[3339] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3340] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'op': 'load'}
    instructions[3341] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3342] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'op': 'load'}
    instructions[3343] = {5'd0, 4'd2, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'literal': 6, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'op': 'literal'}
    instructions[3344] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'op': 'load'}
    instructions[3345] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3346] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'op': 'load'}
    instructions[3347] = {5'd15, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'op': 'not_equal'}
    instructions[3348] = {5'd8, 4'd0, 4'd8, 16'd3361};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'a': 8, 'label': 3361, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'op': 'jmp_if_false'}
    instructions[3349] = {5'd0, 4'd8, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'op': 'literal'}
    instructions[3350] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'op': 'store'}
    instructions[3351] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'op': 'addl'}
    instructions[3352] = {5'd1, 4'd8, 4'd4, 16'd1466};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'a': 4, 'literal': 1466, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'op': 'addl'}
    instructions[3353] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'op': 'addl'}
    instructions[3354] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'op': 'load'}
    instructions[3355] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3356] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'op': 'load'}
    instructions[3357] = {5'd16, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'op': 'or'}
    instructions[3358] = {5'd1, 4'd2, 4'd4, 16'd1466};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'a': 4, 'literal': 1466, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'op': 'addl'}
    instructions[3359] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'op': 'store'}
    instructions[3360] = {5'd12, 4'd0, 4'd0, 16'd3361};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117 {'label': 3361, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 117, 'op': 'goto'}
    instructions[3361] = {5'd0, 4'd8, 4'd0, 16'd65535};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'literal': 65535, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'op': 'literal'}
    instructions[3362] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'op': 'store'}
    instructions[3363] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'op': 'addl'}
    instructions[3364] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'op': 'store'}
    instructions[3365] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'op': 'addl'}
    instructions[3366] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'op': 'store'}
    instructions[3367] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'op': 'addl'}
    instructions[3368] = {5'd1, 4'd8, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'a': 4, 'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'op': 'addl'}
    instructions[3369] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'op': 'store'}
    instructions[3370] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'op': 'addl'}
    instructions[3371] = {5'd0, 4'd8, 4'd0, 16'd67};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'literal': 67, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'op': 'literal'}
    instructions[3372] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'op': 'store'}
    instructions[3373] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'op': 'addl'}
    instructions[3374] = {5'd1, 4'd8, 4'd4, 16'd1467};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'a': 4, 'literal': 1467, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'op': 'addl'}
    instructions[3375] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'op': 'addl'}
    instructions[3376] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'op': 'load'}
    instructions[3377] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'op': 'store'}
    instructions[3378] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'op': 'addl'}
    instructions[3379] = {5'd1, 4'd8, 4'd4, 16'd1468};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'a': 4, 'literal': 1468, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'op': 'addl'}
    instructions[3380] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'op': 'addl'}
    instructions[3381] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'op': 'load'}
    instructions[3382] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'op': 'store'}
    instructions[3383] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'op': 'addl'}
    instructions[3384] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'op': 'addl'}
    instructions[3385] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'op': 'addl'}
    instructions[3386] = {5'd3, 4'd6, 4'd0, 16'd4588};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'z': 6, 'label': 4588, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'op': 'call'}
    instructions[3387] = {5'd1, 4'd3, 4'd3, -16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'a': 3, 'literal': -4, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'op': 'addl'}
    instructions[3388] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3389] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'op': 'load'}
    instructions[3390] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3391] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'op': 'load'}
    instructions[3392] = {5'd0, 4'd2, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'literal': 6, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'op': 'literal'}
    instructions[3393] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'op': 'load'}
    instructions[3394] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3395] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'op': 'load'}
    instructions[3396] = {5'd15, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'op': 'not_equal'}
    instructions[3397] = {5'd8, 4'd0, 4'd8, 16'd3410};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'a': 8, 'label': 3410, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'op': 'jmp_if_false'}
    instructions[3398] = {5'd0, 4'd8, 4'd0, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'literal': 4, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'op': 'literal'}
    instructions[3399] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'op': 'store'}
    instructions[3400] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'op': 'addl'}
    instructions[3401] = {5'd1, 4'd8, 4'd4, 16'd1466};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'a': 4, 'literal': 1466, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'op': 'addl'}
    instructions[3402] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'op': 'addl'}
    instructions[3403] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'op': 'load'}
    instructions[3404] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3405] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'op': 'load'}
    instructions[3406] = {5'd16, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'op': 'or'}
    instructions[3407] = {5'd1, 4'd2, 4'd4, 16'd1466};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'a': 4, 'literal': 1466, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'op': 'addl'}
    instructions[3408] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'op': 'store'}
    instructions[3409] = {5'd12, 4'd0, 4'd0, 16'd3410};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118 {'label': 3410, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 118, 'op': 'goto'}
    instructions[3410] = {5'd0, 4'd8, 4'd0, 16'd65535};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'literal': 65535, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'op': 'literal'}
    instructions[3411] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'op': 'store'}
    instructions[3412] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'op': 'addl'}
    instructions[3413] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'op': 'store'}
    instructions[3414] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'op': 'addl'}
    instructions[3415] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'op': 'store'}
    instructions[3416] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'op': 'addl'}
    instructions[3417] = {5'd1, 4'd8, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'a': 4, 'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'op': 'addl'}
    instructions[3418] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'op': 'store'}
    instructions[3419] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'op': 'addl'}
    instructions[3420] = {5'd0, 4'd8, 4'd0, 16'd68};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'literal': 68, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'op': 'literal'}
    instructions[3421] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'op': 'store'}
    instructions[3422] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'op': 'addl'}
    instructions[3423] = {5'd1, 4'd8, 4'd4, 16'd1467};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'a': 4, 'literal': 1467, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'op': 'addl'}
    instructions[3424] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'op': 'addl'}
    instructions[3425] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'op': 'load'}
    instructions[3426] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'op': 'store'}
    instructions[3427] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'op': 'addl'}
    instructions[3428] = {5'd1, 4'd8, 4'd4, 16'd1468};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'a': 4, 'literal': 1468, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'op': 'addl'}
    instructions[3429] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'op': 'addl'}
    instructions[3430] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'op': 'load'}
    instructions[3431] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'op': 'store'}
    instructions[3432] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'op': 'addl'}
    instructions[3433] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'op': 'addl'}
    instructions[3434] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'op': 'addl'}
    instructions[3435] = {5'd3, 4'd6, 4'd0, 16'd4588};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'z': 6, 'label': 4588, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'op': 'call'}
    instructions[3436] = {5'd1, 4'd3, 4'd3, -16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'a': 3, 'literal': -4, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'op': 'addl'}
    instructions[3437] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3438] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'op': 'load'}
    instructions[3439] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3440] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'op': 'load'}
    instructions[3441] = {5'd0, 4'd2, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'literal': 6, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'op': 'literal'}
    instructions[3442] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'op': 'load'}
    instructions[3443] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3444] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'op': 'load'}
    instructions[3445] = {5'd15, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'op': 'not_equal'}
    instructions[3446] = {5'd8, 4'd0, 4'd8, 16'd3459};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'a': 8, 'label': 3459, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'op': 'jmp_if_false'}
    instructions[3447] = {5'd0, 4'd8, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'literal': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'op': 'literal'}
    instructions[3448] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'op': 'store'}
    instructions[3449] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'op': 'addl'}
    instructions[3450] = {5'd1, 4'd8, 4'd4, 16'd1466};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'a': 4, 'literal': 1466, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'op': 'addl'}
    instructions[3451] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'op': 'addl'}
    instructions[3452] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'op': 'load'}
    instructions[3453] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3454] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'op': 'load'}
    instructions[3455] = {5'd16, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'op': 'or'}
    instructions[3456] = {5'd1, 4'd2, 4'd4, 16'd1466};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'a': 4, 'literal': 1466, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'op': 'addl'}
    instructions[3457] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'op': 'store'}
    instructions[3458] = {5'd12, 4'd0, 4'd0, 16'd3459};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119 {'label': 3459, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 119, 'op': 'goto'}
    instructions[3459] = {5'd0, 4'd8, 4'd0, 16'd65535};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'literal': 65535, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'op': 'literal'}
    instructions[3460] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'op': 'store'}
    instructions[3461] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'op': 'addl'}
    instructions[3462] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'op': 'store'}
    instructions[3463] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'op': 'addl'}
    instructions[3464] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'op': 'store'}
    instructions[3465] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'op': 'addl'}
    instructions[3466] = {5'd1, 4'd8, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'a': 4, 'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'op': 'addl'}
    instructions[3467] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'op': 'store'}
    instructions[3468] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'op': 'addl'}
    instructions[3469] = {5'd0, 4'd8, 4'd0, 16'd69};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'literal': 69, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'op': 'literal'}
    instructions[3470] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'op': 'store'}
    instructions[3471] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'op': 'addl'}
    instructions[3472] = {5'd1, 4'd8, 4'd4, 16'd1467};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'a': 4, 'literal': 1467, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'op': 'addl'}
    instructions[3473] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'op': 'addl'}
    instructions[3474] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'op': 'load'}
    instructions[3475] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'op': 'store'}
    instructions[3476] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'op': 'addl'}
    instructions[3477] = {5'd1, 4'd8, 4'd4, 16'd1468};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'a': 4, 'literal': 1468, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'op': 'addl'}
    instructions[3478] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'op': 'addl'}
    instructions[3479] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'op': 'load'}
    instructions[3480] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'op': 'store'}
    instructions[3481] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'op': 'addl'}
    instructions[3482] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'op': 'addl'}
    instructions[3483] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'op': 'addl'}
    instructions[3484] = {5'd3, 4'd6, 4'd0, 16'd4588};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'z': 6, 'label': 4588, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'op': 'call'}
    instructions[3485] = {5'd1, 4'd3, 4'd3, -16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'a': 3, 'literal': -4, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'op': 'addl'}
    instructions[3486] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3487] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'op': 'load'}
    instructions[3488] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3489] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'op': 'load'}
    instructions[3490] = {5'd0, 4'd2, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'literal': 6, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'op': 'literal'}
    instructions[3491] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'op': 'load'}
    instructions[3492] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3493] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'op': 'load'}
    instructions[3494] = {5'd15, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'op': 'not_equal'}
    instructions[3495] = {5'd8, 4'd0, 4'd8, 16'd3508};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'a': 8, 'label': 3508, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'op': 'jmp_if_false'}
    instructions[3496] = {5'd0, 4'd8, 4'd0, 16'd16};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'literal': 16, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'op': 'literal'}
    instructions[3497] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'op': 'store'}
    instructions[3498] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'op': 'addl'}
    instructions[3499] = {5'd1, 4'd8, 4'd4, 16'd1466};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'a': 4, 'literal': 1466, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'op': 'addl'}
    instructions[3500] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'op': 'addl'}
    instructions[3501] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'op': 'load'}
    instructions[3502] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3503] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'op': 'load'}
    instructions[3504] = {5'd16, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'op': 'or'}
    instructions[3505] = {5'd1, 4'd2, 4'd4, 16'd1466};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'a': 4, 'literal': 1466, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'op': 'addl'}
    instructions[3506] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'op': 'store'}
    instructions[3507] = {5'd12, 4'd0, 4'd0, 16'd3508};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120 {'label': 3508, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 120, 'op': 'goto'}
    instructions[3508] = {5'd0, 4'd8, 4'd0, 16'd65535};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'literal': 65535, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'op': 'literal'}
    instructions[3509] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'op': 'store'}
    instructions[3510] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'op': 'addl'}
    instructions[3511] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'op': 'store'}
    instructions[3512] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'op': 'addl'}
    instructions[3513] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'op': 'store'}
    instructions[3514] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'op': 'addl'}
    instructions[3515] = {5'd1, 4'd8, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'a': 4, 'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'op': 'addl'}
    instructions[3516] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'op': 'store'}
    instructions[3517] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'op': 'addl'}
    instructions[3518] = {5'd0, 4'd8, 4'd0, 16'd70};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'literal': 70, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'op': 'literal'}
    instructions[3519] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'op': 'store'}
    instructions[3520] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'op': 'addl'}
    instructions[3521] = {5'd1, 4'd8, 4'd4, 16'd1467};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'a': 4, 'literal': 1467, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'op': 'addl'}
    instructions[3522] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'op': 'addl'}
    instructions[3523] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'op': 'load'}
    instructions[3524] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'op': 'store'}
    instructions[3525] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'op': 'addl'}
    instructions[3526] = {5'd1, 4'd8, 4'd4, 16'd1468};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'a': 4, 'literal': 1468, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'op': 'addl'}
    instructions[3527] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'op': 'addl'}
    instructions[3528] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'op': 'load'}
    instructions[3529] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'op': 'store'}
    instructions[3530] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'op': 'addl'}
    instructions[3531] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'op': 'addl'}
    instructions[3532] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'op': 'addl'}
    instructions[3533] = {5'd3, 4'd6, 4'd0, 16'd4588};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'z': 6, 'label': 4588, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'op': 'call'}
    instructions[3534] = {5'd1, 4'd3, 4'd3, -16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'a': 3, 'literal': -4, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'op': 'addl'}
    instructions[3535] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3536] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'op': 'load'}
    instructions[3537] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3538] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'op': 'load'}
    instructions[3539] = {5'd0, 4'd2, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'literal': 6, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'op': 'literal'}
    instructions[3540] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'op': 'load'}
    instructions[3541] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3542] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'op': 'load'}
    instructions[3543] = {5'd15, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'op': 'not_equal'}
    instructions[3544] = {5'd8, 4'd0, 4'd8, 16'd3557};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'a': 8, 'label': 3557, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'op': 'jmp_if_false'}
    instructions[3545] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'op': 'literal'}
    instructions[3546] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'op': 'store'}
    instructions[3547] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'op': 'addl'}
    instructions[3548] = {5'd1, 4'd8, 4'd4, 16'd1466};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'a': 4, 'literal': 1466, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'op': 'addl'}
    instructions[3549] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'op': 'addl'}
    instructions[3550] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'op': 'load'}
    instructions[3551] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3552] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'op': 'load'}
    instructions[3553] = {5'd16, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'op': 'or'}
    instructions[3554] = {5'd1, 4'd2, 4'd4, 16'd1466};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'a': 4, 'literal': 1466, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'op': 'addl'}
    instructions[3555] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'op': 'store'}
    instructions[3556] = {5'd12, 4'd0, 4'd0, 16'd3557};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121 {'label': 3557, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 121, 'op': 'goto'}
    instructions[3557] = {5'd0, 4'd8, 4'd0, 16'd65535};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'literal': 65535, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'op': 'literal'}
    instructions[3558] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'op': 'store'}
    instructions[3559] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'op': 'addl'}
    instructions[3560] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'op': 'store'}
    instructions[3561] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'op': 'addl'}
    instructions[3562] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'op': 'store'}
    instructions[3563] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'op': 'addl'}
    instructions[3564] = {5'd1, 4'd8, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'a': 4, 'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'op': 'addl'}
    instructions[3565] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'op': 'store'}
    instructions[3566] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'op': 'addl'}
    instructions[3567] = {5'd0, 4'd8, 4'd0, 16'd71};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'literal': 71, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'op': 'literal'}
    instructions[3568] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'op': 'store'}
    instructions[3569] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'op': 'addl'}
    instructions[3570] = {5'd1, 4'd8, 4'd4, 16'd1467};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'a': 4, 'literal': 1467, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'op': 'addl'}
    instructions[3571] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'op': 'addl'}
    instructions[3572] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'op': 'load'}
    instructions[3573] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'op': 'store'}
    instructions[3574] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'op': 'addl'}
    instructions[3575] = {5'd1, 4'd8, 4'd4, 16'd1468};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'a': 4, 'literal': 1468, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'op': 'addl'}
    instructions[3576] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'op': 'addl'}
    instructions[3577] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'op': 'load'}
    instructions[3578] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'op': 'store'}
    instructions[3579] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'op': 'addl'}
    instructions[3580] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'op': 'addl'}
    instructions[3581] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'op': 'addl'}
    instructions[3582] = {5'd3, 4'd6, 4'd0, 16'd4588};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'z': 6, 'label': 4588, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'op': 'call'}
    instructions[3583] = {5'd1, 4'd3, 4'd3, -16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'a': 3, 'literal': -4, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'op': 'addl'}
    instructions[3584] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3585] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'op': 'load'}
    instructions[3586] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3587] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'op': 'load'}
    instructions[3588] = {5'd0, 4'd2, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'literal': 6, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'op': 'literal'}
    instructions[3589] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'op': 'load'}
    instructions[3590] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3591] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'op': 'load'}
    instructions[3592] = {5'd15, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'op': 'not_equal'}
    instructions[3593] = {5'd8, 4'd0, 4'd8, 16'd3606};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'a': 8, 'label': 3606, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'op': 'jmp_if_false'}
    instructions[3594] = {5'd0, 4'd8, 4'd0, 16'd64};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'literal': 64, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'op': 'literal'}
    instructions[3595] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'op': 'store'}
    instructions[3596] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'op': 'addl'}
    instructions[3597] = {5'd1, 4'd8, 4'd4, 16'd1466};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'a': 4, 'literal': 1466, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'op': 'addl'}
    instructions[3598] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'op': 'addl'}
    instructions[3599] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'op': 'load'}
    instructions[3600] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3601] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'op': 'load'}
    instructions[3602] = {5'd16, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'op': 'or'}
    instructions[3603] = {5'd1, 4'd2, 4'd4, 16'd1466};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'a': 4, 'literal': 1466, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'op': 'addl'}
    instructions[3604] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'op': 'store'}
    instructions[3605] = {5'd12, 4'd0, 4'd0, 16'd3606};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122 {'label': 3606, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 122, 'op': 'goto'}
    instructions[3606] = {5'd0, 4'd8, 4'd0, 16'd65535};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'literal': 65535, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'op': 'literal'}
    instructions[3607] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'op': 'store'}
    instructions[3608] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'op': 'addl'}
    instructions[3609] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'op': 'store'}
    instructions[3610] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'op': 'addl'}
    instructions[3611] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'op': 'store'}
    instructions[3612] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'op': 'addl'}
    instructions[3613] = {5'd1, 4'd8, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'a': 4, 'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'op': 'addl'}
    instructions[3614] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'op': 'store'}
    instructions[3615] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'op': 'addl'}
    instructions[3616] = {5'd0, 4'd8, 4'd0, 16'd72};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'literal': 72, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'op': 'literal'}
    instructions[3617] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'op': 'store'}
    instructions[3618] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'op': 'addl'}
    instructions[3619] = {5'd1, 4'd8, 4'd4, 16'd1467};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'a': 4, 'literal': 1467, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'op': 'addl'}
    instructions[3620] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'op': 'addl'}
    instructions[3621] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'op': 'load'}
    instructions[3622] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'op': 'store'}
    instructions[3623] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'op': 'addl'}
    instructions[3624] = {5'd1, 4'd8, 4'd4, 16'd1468};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'a': 4, 'literal': 1468, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'op': 'addl'}
    instructions[3625] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'op': 'addl'}
    instructions[3626] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'op': 'load'}
    instructions[3627] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'op': 'store'}
    instructions[3628] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'op': 'addl'}
    instructions[3629] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'op': 'addl'}
    instructions[3630] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'op': 'addl'}
    instructions[3631] = {5'd3, 4'd6, 4'd0, 16'd4588};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'z': 6, 'label': 4588, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'op': 'call'}
    instructions[3632] = {5'd1, 4'd3, 4'd3, -16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'a': 3, 'literal': -4, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'op': 'addl'}
    instructions[3633] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3634] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'op': 'load'}
    instructions[3635] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3636] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'op': 'load'}
    instructions[3637] = {5'd0, 4'd2, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'literal': 6, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'op': 'literal'}
    instructions[3638] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'op': 'load'}
    instructions[3639] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3640] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'op': 'load'}
    instructions[3641] = {5'd15, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'op': 'not_equal'}
    instructions[3642] = {5'd8, 4'd0, 4'd8, 16'd3655};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'a': 8, 'label': 3655, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'op': 'jmp_if_false'}
    instructions[3643] = {5'd0, 4'd8, 4'd0, 16'd128};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'literal': 128, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'op': 'literal'}
    instructions[3644] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'op': 'store'}
    instructions[3645] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'op': 'addl'}
    instructions[3646] = {5'd1, 4'd8, 4'd4, 16'd1466};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'a': 4, 'literal': 1466, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'op': 'addl'}
    instructions[3647] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'op': 'addl'}
    instructions[3648] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'op': 'load'}
    instructions[3649] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3650] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'op': 'load'}
    instructions[3651] = {5'd16, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'op': 'or'}
    instructions[3652] = {5'd1, 4'd2, 4'd4, 16'd1466};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'a': 4, 'literal': 1466, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'op': 'addl'}
    instructions[3653] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'op': 'store'}
    instructions[3654] = {5'd12, 4'd0, 4'd0, 16'd3655};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123 {'label': 3655, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 123, 'op': 'goto'}
    instructions[3655] = {5'd0, 4'd8, 4'd0, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 124 {'literal': 10, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 124, 'op': 'literal'}
    instructions[3656] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 124 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 124, 'op': 'addl'}
    instructions[3657] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 124 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 124, 'op': 'load'}
    instructions[3658] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 124 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 124, 'op': 'store'}
    instructions[3659] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 124 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 124, 'op': 'addl'}
    instructions[3660] = {5'd1, 4'd8, 4'd4, 16'd1466};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 124 {'a': 4, 'literal': 1466, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 124, 'op': 'addl'}
    instructions[3661] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 124 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 124, 'op': 'addl'}
    instructions[3662] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 124 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 124, 'op': 'load'}
    instructions[3663] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 124 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 124, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3664] = {5'd5, 4'd0, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 124 {'a': 3, 'z': 0, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 124, 'op': 'load'}
    instructions[3665] = {5'd17, 4'd0, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 124 {'a': 0, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 124, 'op': 'write'}
    instructions[3666] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 124 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 124, 'op': 'addl'}
    instructions[3667] = {5'd0, 4'd8, 4'd0, 16'd11};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 128 {'literal': 11, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 128, 'op': 'literal'}
    instructions[3668] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 128 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 128, 'op': 'addl'}
    instructions[3669] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 128 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 128, 'op': 'load'}
    instructions[3670] = {5'd6, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 128 {'a': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 128, 'op': 'read'}
    instructions[3671] = {5'd18, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 128 {'a': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 128, 'op': 'not'}
    instructions[3672] = {5'd1, 4'd2, 4'd4, 16'd1464};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 128 {'a': 4, 'literal': 1464, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 128, 'op': 'addl'}
    instructions[3673] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 128 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 128, 'op': 'store'}
    instructions[3674] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130, 'op': 'store'}
    instructions[3675] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130, 'op': 'addl'}
    instructions[3676] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130, 'op': 'store'}
    instructions[3677] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130, 'op': 'addl'}
    instructions[3678] = {5'd1, 4'd8, 4'd4, 16'd1469};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130 {'a': 4, 'literal': 1469, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130, 'op': 'addl'}
    instructions[3679] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130, 'op': 'store'}
    instructions[3680] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130, 'op': 'addl'}
    instructions[3681] = {5'd0, 4'd8, 4'd0, 16'd58};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130 {'literal': 58, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130, 'op': 'literal'}
    instructions[3682] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130, 'op': 'store'}
    instructions[3683] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130, 'op': 'addl'}
    instructions[3684] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130, 'op': 'literal'}
    instructions[3685] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130, 'op': 'store'}
    instructions[3686] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130, 'op': 'addl'}
    instructions[3687] = {5'd0, 4'd8, 4'd0, 16'd1460};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130 {'literal': 1460, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130, 'op': 'literal'}
    instructions[3688] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130, 'op': 'store'}
    instructions[3689] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130, 'op': 'addl'}
    instructions[3690] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130, 'op': 'addl'}
    instructions[3691] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130, 'op': 'addl'}
    instructions[3692] = {5'd3, 4'd6, 4'd0, 16'd4588};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130 {'z': 6, 'label': 4588, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130, 'op': 'call'}
    instructions[3693] = {5'd1, 4'd3, 4'd3, -16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130 {'a': 3, 'literal': -4, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130, 'op': 'addl'}
    instructions[3694] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3695] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130, 'op': 'load'}
    instructions[3696] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3697] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130, 'op': 'load'}
    instructions[3698] = {5'd0, 4'd2, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130 {'literal': 6, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130, 'op': 'literal'}
    instructions[3699] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130, 'op': 'load'}
    instructions[3700] = {5'd1, 4'd2, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130 {'a': 4, 'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130, 'op': 'addl'}
    instructions[3701] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 130, 'op': 'store'}
    instructions[3702] = {5'd0, 4'd8, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 131 {'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 131, 'op': 'literal'}
    instructions[3703] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 131 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 131, 'op': 'store'}
    instructions[3704] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 131 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 131, 'op': 'addl'}
    instructions[3705] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 131 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 131, 'op': 'addl'}
    instructions[3706] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 131 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 131, 'op': 'addl'}
    instructions[3707] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 131 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 131, 'op': 'load'}
    instructions[3708] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 131 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 131, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3709] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 131 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 131, 'op': 'load'}
    instructions[3710] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 131 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 131, 'op': 'add'}
    instructions[3711] = {5'd1, 4'd2, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 131 {'a': 4, 'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 131, 'op': 'addl'}
    instructions[3712] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 131 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 131, 'op': 'store'}
    instructions[3713] = {5'd0, 4'd8, 4'd0, 16'd128};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133 {'literal': 128, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133, 'op': 'literal'}
    instructions[3714] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133, 'op': 'store'}
    instructions[3715] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133, 'op': 'addl'}
    instructions[3716] = {5'd1, 4'd8, 4'd4, 16'd1464};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133 {'a': 4, 'literal': 1464, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133, 'op': 'addl'}
    instructions[3717] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133, 'op': 'addl'}
    instructions[3718] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133, 'op': 'load'}
    instructions[3719] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3720] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133, 'op': 'load'}
    instructions[3721] = {5'd10, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133, 'op': 'and'}
    instructions[3722] = {5'd8, 4'd0, 4'd8, 16'd3740};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133 {'a': 8, 'label': 3740, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133, 'op': 'jmp_if_false'}
    instructions[3723] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133, 'op': 'literal'}
    instructions[3724] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133, 'op': 'store'}
    instructions[3725] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133, 'op': 'addl'}
    instructions[3726] = {5'd1, 4'd8, 4'd4, 16'd1469};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133 {'a': 4, 'literal': 1469, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133, 'op': 'addl'}
    instructions[3727] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133, 'op': 'store'}
    instructions[3728] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133, 'op': 'addl'}
    instructions[3729] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133, 'op': 'addl'}
    instructions[3730] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133, 'op': 'addl'}
    instructions[3731] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133, 'op': 'load'}
    instructions[3732] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3733] = {5'd5, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133, 'op': 'load'}
    instructions[3734] = {5'd11, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133, 'op': 'add'}
    instructions[3735] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133, 'op': 'addl'}
    instructions[3736] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3737] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133, 'op': 'load'}
    instructions[3738] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133, 'op': 'store'}
    instructions[3739] = {5'd12, 4'd0, 4'd0, 16'd3756};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133 {'label': 3756, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 133, 'op': 'goto'}
    instructions[3740] = {5'd0, 4'd8, 4'd0, 16'd49};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 134 {'literal': 49, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 134, 'op': 'literal'}
    instructions[3741] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 134 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 134, 'op': 'store'}
    instructions[3742] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 134 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 134, 'op': 'addl'}
    instructions[3743] = {5'd1, 4'd8, 4'd4, 16'd1469};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 134 {'a': 4, 'literal': 1469, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 134, 'op': 'addl'}
    instructions[3744] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 134 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 134, 'op': 'store'}
    instructions[3745] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 134 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 134, 'op': 'addl'}
    instructions[3746] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 134 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 134, 'op': 'addl'}
    instructions[3747] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 134 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 134, 'op': 'addl'}
    instructions[3748] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 134 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 134, 'op': 'load'}
    instructions[3749] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 134 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 134, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3750] = {5'd5, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 134 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 134, 'op': 'load'}
    instructions[3751] = {5'd11, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 134 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 134, 'op': 'add'}
    instructions[3752] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 134 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 134, 'op': 'addl'}
    instructions[3753] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 134 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 134, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3754] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 134 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 134, 'op': 'load'}
    instructions[3755] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 134 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 134, 'op': 'store'}
    instructions[3756] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 135 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 135, 'op': 'addl'}
    instructions[3757] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 135 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 135, 'op': 'addl'}
    instructions[3758] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 135 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 135, 'op': 'load'}
    instructions[3759] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 135 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 135, 'op': 'store'}
    instructions[3760] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 135 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 135, 'op': 'addl'}
    instructions[3761] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 135 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 135, 'op': 'literal'}
    instructions[3762] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 135 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 135, 'op': 'store'}
    instructions[3763] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 135 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 135, 'op': 'addl'}
    instructions[3764] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 135 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 135, 'op': 'addl'}
    instructions[3765] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 135 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 135, 'op': 'addl'}
    instructions[3766] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 135 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 135, 'op': 'load'}
    instructions[3767] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 135 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 135, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3768] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 135 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 135, 'op': 'load'}
    instructions[3769] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 135 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 135, 'op': 'add'}
    instructions[3770] = {5'd1, 4'd2, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 135 {'a': 4, 'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 135, 'op': 'addl'}
    instructions[3771] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 135 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 135, 'op': 'store'}
    instructions[3772] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 135 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 135, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3773] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 135 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 135, 'op': 'load'}
    instructions[3774] = {5'd0, 4'd8, 4'd0, 16'd64};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136 {'literal': 64, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136, 'op': 'literal'}
    instructions[3775] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136, 'op': 'store'}
    instructions[3776] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136, 'op': 'addl'}
    instructions[3777] = {5'd1, 4'd8, 4'd4, 16'd1464};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136 {'a': 4, 'literal': 1464, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136, 'op': 'addl'}
    instructions[3778] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136, 'op': 'addl'}
    instructions[3779] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136, 'op': 'load'}
    instructions[3780] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3781] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136, 'op': 'load'}
    instructions[3782] = {5'd10, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136, 'op': 'and'}
    instructions[3783] = {5'd8, 4'd0, 4'd8, 16'd3801};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136 {'a': 8, 'label': 3801, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136, 'op': 'jmp_if_false'}
    instructions[3784] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136, 'op': 'literal'}
    instructions[3785] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136, 'op': 'store'}
    instructions[3786] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136, 'op': 'addl'}
    instructions[3787] = {5'd1, 4'd8, 4'd4, 16'd1469};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136 {'a': 4, 'literal': 1469, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136, 'op': 'addl'}
    instructions[3788] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136, 'op': 'store'}
    instructions[3789] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136, 'op': 'addl'}
    instructions[3790] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136, 'op': 'addl'}
    instructions[3791] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136, 'op': 'addl'}
    instructions[3792] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136, 'op': 'load'}
    instructions[3793] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3794] = {5'd5, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136, 'op': 'load'}
    instructions[3795] = {5'd11, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136, 'op': 'add'}
    instructions[3796] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136, 'op': 'addl'}
    instructions[3797] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3798] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136, 'op': 'load'}
    instructions[3799] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136, 'op': 'store'}
    instructions[3800] = {5'd12, 4'd0, 4'd0, 16'd3817};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136 {'label': 3817, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 136, 'op': 'goto'}
    instructions[3801] = {5'd0, 4'd8, 4'd0, 16'd49};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 137 {'literal': 49, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 137, 'op': 'literal'}
    instructions[3802] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 137 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 137, 'op': 'store'}
    instructions[3803] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 137 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 137, 'op': 'addl'}
    instructions[3804] = {5'd1, 4'd8, 4'd4, 16'd1469};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 137 {'a': 4, 'literal': 1469, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 137, 'op': 'addl'}
    instructions[3805] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 137 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 137, 'op': 'store'}
    instructions[3806] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 137 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 137, 'op': 'addl'}
    instructions[3807] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 137 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 137, 'op': 'addl'}
    instructions[3808] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 137 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 137, 'op': 'addl'}
    instructions[3809] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 137 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 137, 'op': 'load'}
    instructions[3810] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 137 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 137, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3811] = {5'd5, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 137 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 137, 'op': 'load'}
    instructions[3812] = {5'd11, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 137 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 137, 'op': 'add'}
    instructions[3813] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 137 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 137, 'op': 'addl'}
    instructions[3814] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 137 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 137, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3815] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 137 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 137, 'op': 'load'}
    instructions[3816] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 137 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 137, 'op': 'store'}
    instructions[3817] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 138 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 138, 'op': 'addl'}
    instructions[3818] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 138 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 138, 'op': 'addl'}
    instructions[3819] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 138 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 138, 'op': 'load'}
    instructions[3820] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 138 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 138, 'op': 'store'}
    instructions[3821] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 138 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 138, 'op': 'addl'}
    instructions[3822] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 138 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 138, 'op': 'literal'}
    instructions[3823] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 138 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 138, 'op': 'store'}
    instructions[3824] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 138 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 138, 'op': 'addl'}
    instructions[3825] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 138 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 138, 'op': 'addl'}
    instructions[3826] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 138 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 138, 'op': 'addl'}
    instructions[3827] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 138 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 138, 'op': 'load'}
    instructions[3828] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 138 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 138, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3829] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 138 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 138, 'op': 'load'}
    instructions[3830] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 138 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 138, 'op': 'add'}
    instructions[3831] = {5'd1, 4'd2, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 138 {'a': 4, 'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 138, 'op': 'addl'}
    instructions[3832] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 138 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 138, 'op': 'store'}
    instructions[3833] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 138 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 138, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3834] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 138 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 138, 'op': 'load'}
    instructions[3835] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139, 'op': 'literal'}
    instructions[3836] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139, 'op': 'store'}
    instructions[3837] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139, 'op': 'addl'}
    instructions[3838] = {5'd1, 4'd8, 4'd4, 16'd1464};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139 {'a': 4, 'literal': 1464, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139, 'op': 'addl'}
    instructions[3839] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139, 'op': 'addl'}
    instructions[3840] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139, 'op': 'load'}
    instructions[3841] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3842] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139, 'op': 'load'}
    instructions[3843] = {5'd10, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139, 'op': 'and'}
    instructions[3844] = {5'd8, 4'd0, 4'd8, 16'd3862};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139 {'a': 8, 'label': 3862, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139, 'op': 'jmp_if_false'}
    instructions[3845] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139, 'op': 'literal'}
    instructions[3846] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139, 'op': 'store'}
    instructions[3847] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139, 'op': 'addl'}
    instructions[3848] = {5'd1, 4'd8, 4'd4, 16'd1469};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139 {'a': 4, 'literal': 1469, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139, 'op': 'addl'}
    instructions[3849] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139, 'op': 'store'}
    instructions[3850] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139, 'op': 'addl'}
    instructions[3851] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139, 'op': 'addl'}
    instructions[3852] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139, 'op': 'addl'}
    instructions[3853] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139, 'op': 'load'}
    instructions[3854] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3855] = {5'd5, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139, 'op': 'load'}
    instructions[3856] = {5'd11, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139, 'op': 'add'}
    instructions[3857] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139, 'op': 'addl'}
    instructions[3858] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3859] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139, 'op': 'load'}
    instructions[3860] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139, 'op': 'store'}
    instructions[3861] = {5'd12, 4'd0, 4'd0, 16'd3878};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139 {'label': 3878, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 139, 'op': 'goto'}
    instructions[3862] = {5'd0, 4'd8, 4'd0, 16'd49};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 140 {'literal': 49, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 140, 'op': 'literal'}
    instructions[3863] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 140 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 140, 'op': 'store'}
    instructions[3864] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 140 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 140, 'op': 'addl'}
    instructions[3865] = {5'd1, 4'd8, 4'd4, 16'd1469};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 140 {'a': 4, 'literal': 1469, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 140, 'op': 'addl'}
    instructions[3866] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 140 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 140, 'op': 'store'}
    instructions[3867] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 140 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 140, 'op': 'addl'}
    instructions[3868] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 140 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 140, 'op': 'addl'}
    instructions[3869] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 140 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 140, 'op': 'addl'}
    instructions[3870] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 140 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 140, 'op': 'load'}
    instructions[3871] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 140 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 140, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3872] = {5'd5, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 140 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 140, 'op': 'load'}
    instructions[3873] = {5'd11, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 140 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 140, 'op': 'add'}
    instructions[3874] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 140 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 140, 'op': 'addl'}
    instructions[3875] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 140 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 140, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3876] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 140 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 140, 'op': 'load'}
    instructions[3877] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 140 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 140, 'op': 'store'}
    instructions[3878] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 141 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 141, 'op': 'addl'}
    instructions[3879] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 141 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 141, 'op': 'addl'}
    instructions[3880] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 141 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 141, 'op': 'load'}
    instructions[3881] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 141 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 141, 'op': 'store'}
    instructions[3882] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 141 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 141, 'op': 'addl'}
    instructions[3883] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 141 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 141, 'op': 'literal'}
    instructions[3884] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 141 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 141, 'op': 'store'}
    instructions[3885] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 141 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 141, 'op': 'addl'}
    instructions[3886] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 141 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 141, 'op': 'addl'}
    instructions[3887] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 141 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 141, 'op': 'addl'}
    instructions[3888] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 141 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 141, 'op': 'load'}
    instructions[3889] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 141 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 141, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3890] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 141 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 141, 'op': 'load'}
    instructions[3891] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 141 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 141, 'op': 'add'}
    instructions[3892] = {5'd1, 4'd2, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 141 {'a': 4, 'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 141, 'op': 'addl'}
    instructions[3893] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 141 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 141, 'op': 'store'}
    instructions[3894] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 141 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 141, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3895] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 141 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 141, 'op': 'load'}
    instructions[3896] = {5'd0, 4'd8, 4'd0, 16'd16};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142 {'literal': 16, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142, 'op': 'literal'}
    instructions[3897] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142, 'op': 'store'}
    instructions[3898] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142, 'op': 'addl'}
    instructions[3899] = {5'd1, 4'd8, 4'd4, 16'd1464};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142 {'a': 4, 'literal': 1464, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142, 'op': 'addl'}
    instructions[3900] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142, 'op': 'addl'}
    instructions[3901] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142, 'op': 'load'}
    instructions[3902] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3903] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142, 'op': 'load'}
    instructions[3904] = {5'd10, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142, 'op': 'and'}
    instructions[3905] = {5'd8, 4'd0, 4'd8, 16'd3923};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142 {'a': 8, 'label': 3923, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142, 'op': 'jmp_if_false'}
    instructions[3906] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142, 'op': 'literal'}
    instructions[3907] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142, 'op': 'store'}
    instructions[3908] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142, 'op': 'addl'}
    instructions[3909] = {5'd1, 4'd8, 4'd4, 16'd1469};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142 {'a': 4, 'literal': 1469, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142, 'op': 'addl'}
    instructions[3910] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142, 'op': 'store'}
    instructions[3911] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142, 'op': 'addl'}
    instructions[3912] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142, 'op': 'addl'}
    instructions[3913] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142, 'op': 'addl'}
    instructions[3914] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142, 'op': 'load'}
    instructions[3915] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3916] = {5'd5, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142, 'op': 'load'}
    instructions[3917] = {5'd11, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142, 'op': 'add'}
    instructions[3918] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142, 'op': 'addl'}
    instructions[3919] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3920] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142, 'op': 'load'}
    instructions[3921] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142, 'op': 'store'}
    instructions[3922] = {5'd12, 4'd0, 4'd0, 16'd3939};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142 {'label': 3939, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 142, 'op': 'goto'}
    instructions[3923] = {5'd0, 4'd8, 4'd0, 16'd49};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 143 {'literal': 49, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 143, 'op': 'literal'}
    instructions[3924] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 143 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 143, 'op': 'store'}
    instructions[3925] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 143 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 143, 'op': 'addl'}
    instructions[3926] = {5'd1, 4'd8, 4'd4, 16'd1469};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 143 {'a': 4, 'literal': 1469, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 143, 'op': 'addl'}
    instructions[3927] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 143 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 143, 'op': 'store'}
    instructions[3928] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 143 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 143, 'op': 'addl'}
    instructions[3929] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 143 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 143, 'op': 'addl'}
    instructions[3930] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 143 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 143, 'op': 'addl'}
    instructions[3931] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 143 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 143, 'op': 'load'}
    instructions[3932] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 143 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 143, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3933] = {5'd5, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 143 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 143, 'op': 'load'}
    instructions[3934] = {5'd11, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 143 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 143, 'op': 'add'}
    instructions[3935] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 143 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 143, 'op': 'addl'}
    instructions[3936] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 143 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 143, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3937] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 143 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 143, 'op': 'load'}
    instructions[3938] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 143 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 143, 'op': 'store'}
    instructions[3939] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 144 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 144, 'op': 'addl'}
    instructions[3940] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 144 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 144, 'op': 'addl'}
    instructions[3941] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 144 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 144, 'op': 'load'}
    instructions[3942] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 144 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 144, 'op': 'store'}
    instructions[3943] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 144 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 144, 'op': 'addl'}
    instructions[3944] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 144 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 144, 'op': 'literal'}
    instructions[3945] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 144 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 144, 'op': 'store'}
    instructions[3946] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 144 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 144, 'op': 'addl'}
    instructions[3947] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 144 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 144, 'op': 'addl'}
    instructions[3948] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 144 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 144, 'op': 'addl'}
    instructions[3949] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 144 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 144, 'op': 'load'}
    instructions[3950] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 144 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 144, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3951] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 144 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 144, 'op': 'load'}
    instructions[3952] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 144 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 144, 'op': 'add'}
    instructions[3953] = {5'd1, 4'd2, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 144 {'a': 4, 'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 144, 'op': 'addl'}
    instructions[3954] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 144 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 144, 'op': 'store'}
    instructions[3955] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 144 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 144, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3956] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 144 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 144, 'op': 'load'}
    instructions[3957] = {5'd0, 4'd8, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145 {'literal': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145, 'op': 'literal'}
    instructions[3958] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145, 'op': 'store'}
    instructions[3959] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145, 'op': 'addl'}
    instructions[3960] = {5'd1, 4'd8, 4'd4, 16'd1464};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145 {'a': 4, 'literal': 1464, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145, 'op': 'addl'}
    instructions[3961] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145, 'op': 'addl'}
    instructions[3962] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145, 'op': 'load'}
    instructions[3963] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3964] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145, 'op': 'load'}
    instructions[3965] = {5'd10, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145, 'op': 'and'}
    instructions[3966] = {5'd8, 4'd0, 4'd8, 16'd3984};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145 {'a': 8, 'label': 3984, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145, 'op': 'jmp_if_false'}
    instructions[3967] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145, 'op': 'literal'}
    instructions[3968] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145, 'op': 'store'}
    instructions[3969] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145, 'op': 'addl'}
    instructions[3970] = {5'd1, 4'd8, 4'd4, 16'd1469};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145 {'a': 4, 'literal': 1469, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145, 'op': 'addl'}
    instructions[3971] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145, 'op': 'store'}
    instructions[3972] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145, 'op': 'addl'}
    instructions[3973] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145, 'op': 'addl'}
    instructions[3974] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145, 'op': 'addl'}
    instructions[3975] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145, 'op': 'load'}
    instructions[3976] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3977] = {5'd5, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145, 'op': 'load'}
    instructions[3978] = {5'd11, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145, 'op': 'add'}
    instructions[3979] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145, 'op': 'addl'}
    instructions[3980] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3981] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145, 'op': 'load'}
    instructions[3982] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145, 'op': 'store'}
    instructions[3983] = {5'd12, 4'd0, 4'd0, 16'd4000};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145 {'label': 4000, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 145, 'op': 'goto'}
    instructions[3984] = {5'd0, 4'd8, 4'd0, 16'd49};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 146 {'literal': 49, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 146, 'op': 'literal'}
    instructions[3985] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 146 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 146, 'op': 'store'}
    instructions[3986] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 146 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 146, 'op': 'addl'}
    instructions[3987] = {5'd1, 4'd8, 4'd4, 16'd1469};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 146 {'a': 4, 'literal': 1469, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 146, 'op': 'addl'}
    instructions[3988] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 146 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 146, 'op': 'store'}
    instructions[3989] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 146 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 146, 'op': 'addl'}
    instructions[3990] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 146 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 146, 'op': 'addl'}
    instructions[3991] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 146 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 146, 'op': 'addl'}
    instructions[3992] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 146 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 146, 'op': 'load'}
    instructions[3993] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 146 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 146, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3994] = {5'd5, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 146 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 146, 'op': 'load'}
    instructions[3995] = {5'd11, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 146 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 146, 'op': 'add'}
    instructions[3996] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 146 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 146, 'op': 'addl'}
    instructions[3997] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 146 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 146, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3998] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 146 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 146, 'op': 'load'}
    instructions[3999] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 146 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 146, 'op': 'store'}
    instructions[4000] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 147 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 147, 'op': 'addl'}
    instructions[4001] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 147 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 147, 'op': 'addl'}
    instructions[4002] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 147 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 147, 'op': 'load'}
    instructions[4003] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 147 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 147, 'op': 'store'}
    instructions[4004] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 147 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 147, 'op': 'addl'}
    instructions[4005] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 147 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 147, 'op': 'literal'}
    instructions[4006] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 147 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 147, 'op': 'store'}
    instructions[4007] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 147 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 147, 'op': 'addl'}
    instructions[4008] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 147 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 147, 'op': 'addl'}
    instructions[4009] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 147 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 147, 'op': 'addl'}
    instructions[4010] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 147 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 147, 'op': 'load'}
    instructions[4011] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 147 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 147, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4012] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 147 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 147, 'op': 'load'}
    instructions[4013] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 147 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 147, 'op': 'add'}
    instructions[4014] = {5'd1, 4'd2, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 147 {'a': 4, 'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 147, 'op': 'addl'}
    instructions[4015] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 147 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 147, 'op': 'store'}
    instructions[4016] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 147 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 147, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4017] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 147 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 147, 'op': 'load'}
    instructions[4018] = {5'd0, 4'd8, 4'd0, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148 {'literal': 4, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148, 'op': 'literal'}
    instructions[4019] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148, 'op': 'store'}
    instructions[4020] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148, 'op': 'addl'}
    instructions[4021] = {5'd1, 4'd8, 4'd4, 16'd1464};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148 {'a': 4, 'literal': 1464, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148, 'op': 'addl'}
    instructions[4022] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148, 'op': 'addl'}
    instructions[4023] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148, 'op': 'load'}
    instructions[4024] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4025] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148, 'op': 'load'}
    instructions[4026] = {5'd10, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148, 'op': 'and'}
    instructions[4027] = {5'd8, 4'd0, 4'd8, 16'd4045};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148 {'a': 8, 'label': 4045, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148, 'op': 'jmp_if_false'}
    instructions[4028] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148, 'op': 'literal'}
    instructions[4029] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148, 'op': 'store'}
    instructions[4030] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148, 'op': 'addl'}
    instructions[4031] = {5'd1, 4'd8, 4'd4, 16'd1469};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148 {'a': 4, 'literal': 1469, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148, 'op': 'addl'}
    instructions[4032] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148, 'op': 'store'}
    instructions[4033] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148, 'op': 'addl'}
    instructions[4034] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148, 'op': 'addl'}
    instructions[4035] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148, 'op': 'addl'}
    instructions[4036] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148, 'op': 'load'}
    instructions[4037] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4038] = {5'd5, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148, 'op': 'load'}
    instructions[4039] = {5'd11, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148, 'op': 'add'}
    instructions[4040] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148, 'op': 'addl'}
    instructions[4041] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4042] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148, 'op': 'load'}
    instructions[4043] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148, 'op': 'store'}
    instructions[4044] = {5'd12, 4'd0, 4'd0, 16'd4061};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148 {'label': 4061, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 148, 'op': 'goto'}
    instructions[4045] = {5'd0, 4'd8, 4'd0, 16'd49};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 149 {'literal': 49, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 149, 'op': 'literal'}
    instructions[4046] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 149 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 149, 'op': 'store'}
    instructions[4047] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 149 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 149, 'op': 'addl'}
    instructions[4048] = {5'd1, 4'd8, 4'd4, 16'd1469};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 149 {'a': 4, 'literal': 1469, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 149, 'op': 'addl'}
    instructions[4049] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 149 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 149, 'op': 'store'}
    instructions[4050] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 149 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 149, 'op': 'addl'}
    instructions[4051] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 149 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 149, 'op': 'addl'}
    instructions[4052] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 149 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 149, 'op': 'addl'}
    instructions[4053] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 149 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 149, 'op': 'load'}
    instructions[4054] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 149 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 149, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4055] = {5'd5, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 149 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 149, 'op': 'load'}
    instructions[4056] = {5'd11, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 149 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 149, 'op': 'add'}
    instructions[4057] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 149 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 149, 'op': 'addl'}
    instructions[4058] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 149 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 149, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4059] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 149 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 149, 'op': 'load'}
    instructions[4060] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 149 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 149, 'op': 'store'}
    instructions[4061] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 150 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 150, 'op': 'addl'}
    instructions[4062] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 150 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 150, 'op': 'addl'}
    instructions[4063] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 150 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 150, 'op': 'load'}
    instructions[4064] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 150 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 150, 'op': 'store'}
    instructions[4065] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 150 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 150, 'op': 'addl'}
    instructions[4066] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 150 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 150, 'op': 'literal'}
    instructions[4067] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 150 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 150, 'op': 'store'}
    instructions[4068] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 150 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 150, 'op': 'addl'}
    instructions[4069] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 150 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 150, 'op': 'addl'}
    instructions[4070] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 150 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 150, 'op': 'addl'}
    instructions[4071] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 150 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 150, 'op': 'load'}
    instructions[4072] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 150 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 150, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4073] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 150 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 150, 'op': 'load'}
    instructions[4074] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 150 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 150, 'op': 'add'}
    instructions[4075] = {5'd1, 4'd2, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 150 {'a': 4, 'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 150, 'op': 'addl'}
    instructions[4076] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 150 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 150, 'op': 'store'}
    instructions[4077] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 150 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 150, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4078] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 150 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 150, 'op': 'load'}
    instructions[4079] = {5'd0, 4'd8, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151 {'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151, 'op': 'literal'}
    instructions[4080] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151, 'op': 'store'}
    instructions[4081] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151, 'op': 'addl'}
    instructions[4082] = {5'd1, 4'd8, 4'd4, 16'd1464};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151 {'a': 4, 'literal': 1464, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151, 'op': 'addl'}
    instructions[4083] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151, 'op': 'addl'}
    instructions[4084] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151, 'op': 'load'}
    instructions[4085] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4086] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151, 'op': 'load'}
    instructions[4087] = {5'd10, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151, 'op': 'and'}
    instructions[4088] = {5'd8, 4'd0, 4'd8, 16'd4106};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151 {'a': 8, 'label': 4106, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151, 'op': 'jmp_if_false'}
    instructions[4089] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151, 'op': 'literal'}
    instructions[4090] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151, 'op': 'store'}
    instructions[4091] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151, 'op': 'addl'}
    instructions[4092] = {5'd1, 4'd8, 4'd4, 16'd1469};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151 {'a': 4, 'literal': 1469, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151, 'op': 'addl'}
    instructions[4093] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151, 'op': 'store'}
    instructions[4094] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151, 'op': 'addl'}
    instructions[4095] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151, 'op': 'addl'}
    instructions[4096] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151, 'op': 'addl'}
    instructions[4097] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151, 'op': 'load'}
    instructions[4098] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4099] = {5'd5, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151, 'op': 'load'}
    instructions[4100] = {5'd11, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151, 'op': 'add'}
    instructions[4101] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151, 'op': 'addl'}
    instructions[4102] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4103] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151, 'op': 'load'}
    instructions[4104] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151, 'op': 'store'}
    instructions[4105] = {5'd12, 4'd0, 4'd0, 16'd4122};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151 {'label': 4122, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 151, 'op': 'goto'}
    instructions[4106] = {5'd0, 4'd8, 4'd0, 16'd49};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 152 {'literal': 49, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 152, 'op': 'literal'}
    instructions[4107] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 152 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 152, 'op': 'store'}
    instructions[4108] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 152 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 152, 'op': 'addl'}
    instructions[4109] = {5'd1, 4'd8, 4'd4, 16'd1469};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 152 {'a': 4, 'literal': 1469, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 152, 'op': 'addl'}
    instructions[4110] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 152 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 152, 'op': 'store'}
    instructions[4111] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 152 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 152, 'op': 'addl'}
    instructions[4112] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 152 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 152, 'op': 'addl'}
    instructions[4113] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 152 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 152, 'op': 'addl'}
    instructions[4114] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 152 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 152, 'op': 'load'}
    instructions[4115] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 152 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 152, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4116] = {5'd5, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 152 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 152, 'op': 'load'}
    instructions[4117] = {5'd11, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 152 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 152, 'op': 'add'}
    instructions[4118] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 152 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 152, 'op': 'addl'}
    instructions[4119] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 152 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 152, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4120] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 152 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 152, 'op': 'load'}
    instructions[4121] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 152 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 152, 'op': 'store'}
    instructions[4122] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 153 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 153, 'op': 'addl'}
    instructions[4123] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 153 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 153, 'op': 'addl'}
    instructions[4124] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 153 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 153, 'op': 'load'}
    instructions[4125] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 153 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 153, 'op': 'store'}
    instructions[4126] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 153 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 153, 'op': 'addl'}
    instructions[4127] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 153 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 153, 'op': 'literal'}
    instructions[4128] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 153 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 153, 'op': 'store'}
    instructions[4129] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 153 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 153, 'op': 'addl'}
    instructions[4130] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 153 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 153, 'op': 'addl'}
    instructions[4131] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 153 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 153, 'op': 'addl'}
    instructions[4132] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 153 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 153, 'op': 'load'}
    instructions[4133] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 153 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 153, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4134] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 153 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 153, 'op': 'load'}
    instructions[4135] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 153 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 153, 'op': 'add'}
    instructions[4136] = {5'd1, 4'd2, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 153 {'a': 4, 'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 153, 'op': 'addl'}
    instructions[4137] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 153 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 153, 'op': 'store'}
    instructions[4138] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 153 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 153, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4139] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 153 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 153, 'op': 'load'}
    instructions[4140] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154, 'op': 'literal'}
    instructions[4141] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154, 'op': 'store'}
    instructions[4142] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154, 'op': 'addl'}
    instructions[4143] = {5'd1, 4'd8, 4'd4, 16'd1464};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154 {'a': 4, 'literal': 1464, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154, 'op': 'addl'}
    instructions[4144] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154, 'op': 'addl'}
    instructions[4145] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154, 'op': 'load'}
    instructions[4146] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4147] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154, 'op': 'load'}
    instructions[4148] = {5'd10, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154, 'op': 'and'}
    instructions[4149] = {5'd8, 4'd0, 4'd8, 16'd4167};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154 {'a': 8, 'label': 4167, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154, 'op': 'jmp_if_false'}
    instructions[4150] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154, 'op': 'literal'}
    instructions[4151] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154, 'op': 'store'}
    instructions[4152] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154, 'op': 'addl'}
    instructions[4153] = {5'd1, 4'd8, 4'd4, 16'd1469};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154 {'a': 4, 'literal': 1469, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154, 'op': 'addl'}
    instructions[4154] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154, 'op': 'store'}
    instructions[4155] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154, 'op': 'addl'}
    instructions[4156] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154, 'op': 'addl'}
    instructions[4157] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154, 'op': 'addl'}
    instructions[4158] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154, 'op': 'load'}
    instructions[4159] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4160] = {5'd5, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154, 'op': 'load'}
    instructions[4161] = {5'd11, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154, 'op': 'add'}
    instructions[4162] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154, 'op': 'addl'}
    instructions[4163] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4164] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154, 'op': 'load'}
    instructions[4165] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154, 'op': 'store'}
    instructions[4166] = {5'd12, 4'd0, 4'd0, 16'd4183};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154 {'label': 4183, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 154, 'op': 'goto'}
    instructions[4167] = {5'd0, 4'd8, 4'd0, 16'd49};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 155 {'literal': 49, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 155, 'op': 'literal'}
    instructions[4168] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 155 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 155, 'op': 'store'}
    instructions[4169] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 155 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 155, 'op': 'addl'}
    instructions[4170] = {5'd1, 4'd8, 4'd4, 16'd1469};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 155 {'a': 4, 'literal': 1469, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 155, 'op': 'addl'}
    instructions[4171] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 155 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 155, 'op': 'store'}
    instructions[4172] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 155 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 155, 'op': 'addl'}
    instructions[4173] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 155 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 155, 'op': 'addl'}
    instructions[4174] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 155 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 155, 'op': 'addl'}
    instructions[4175] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 155 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 155, 'op': 'load'}
    instructions[4176] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 155 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 155, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4177] = {5'd5, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 155 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 155, 'op': 'load'}
    instructions[4178] = {5'd11, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 155 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 155, 'op': 'add'}
    instructions[4179] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 155 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 155, 'op': 'addl'}
    instructions[4180] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 155 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 155, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4181] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 155 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 155, 'op': 'load'}
    instructions[4182] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 155 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 155, 'op': 'store'}
    instructions[4183] = {5'd0, 4'd8, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 159 {'literal': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 159, 'op': 'literal'}
    instructions[4184] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 159 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 159, 'op': 'addl'}
    instructions[4185] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 159 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 159, 'op': 'load'}
    instructions[4186] = {5'd6, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 159 {'a': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 159, 'op': 'read'}
    instructions[4187] = {5'd18, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 159 {'a': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 159, 'op': 'not'}
    instructions[4188] = {5'd1, 4'd2, 4'd4, 16'd1465};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 159 {'a': 4, 'literal': 1465, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 159, 'op': 'addl'}
    instructions[4189] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 159 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 159, 'op': 'store'}
    instructions[4190] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161, 'op': 'store'}
    instructions[4191] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161, 'op': 'addl'}
    instructions[4192] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161, 'op': 'store'}
    instructions[4193] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161, 'op': 'addl'}
    instructions[4194] = {5'd1, 4'd8, 4'd4, 16'd1469};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161 {'a': 4, 'literal': 1469, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161, 'op': 'addl'}
    instructions[4195] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161, 'op': 'store'}
    instructions[4196] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161, 'op': 'addl'}
    instructions[4197] = {5'd0, 4'd8, 4'd0, 16'd58};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161 {'literal': 58, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161, 'op': 'literal'}
    instructions[4198] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161, 'op': 'store'}
    instructions[4199] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161, 'op': 'addl'}
    instructions[4200] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161, 'op': 'literal'}
    instructions[4201] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161, 'op': 'store'}
    instructions[4202] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161, 'op': 'addl'}
    instructions[4203] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161, 'op': 'addl'}
    instructions[4204] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161, 'op': 'addl'}
    instructions[4205] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161, 'op': 'load'}
    instructions[4206] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4207] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161, 'op': 'load'}
    instructions[4208] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161, 'op': 'add'}
    instructions[4209] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161, 'op': 'store'}
    instructions[4210] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161, 'op': 'addl'}
    instructions[4211] = {5'd0, 4'd8, 4'd0, 16'd1460};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161 {'literal': 1460, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161, 'op': 'literal'}
    instructions[4212] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161, 'op': 'store'}
    instructions[4213] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161, 'op': 'addl'}
    instructions[4214] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161, 'op': 'addl'}
    instructions[4215] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161, 'op': 'addl'}
    instructions[4216] = {5'd3, 4'd6, 4'd0, 16'd4588};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161 {'z': 6, 'label': 4588, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161, 'op': 'call'}
    instructions[4217] = {5'd1, 4'd3, 4'd3, -16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161 {'a': 3, 'literal': -4, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161, 'op': 'addl'}
    instructions[4218] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4219] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161, 'op': 'load'}
    instructions[4220] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4221] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161, 'op': 'load'}
    instructions[4222] = {5'd0, 4'd2, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161 {'literal': 6, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161, 'op': 'literal'}
    instructions[4223] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161, 'op': 'load'}
    instructions[4224] = {5'd1, 4'd2, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161 {'a': 4, 'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161, 'op': 'addl'}
    instructions[4225] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 161, 'op': 'store'}
    instructions[4226] = {5'd0, 4'd8, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 162 {'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 162, 'op': 'literal'}
    instructions[4227] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 162 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 162, 'op': 'store'}
    instructions[4228] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 162 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 162, 'op': 'addl'}
    instructions[4229] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 162 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 162, 'op': 'addl'}
    instructions[4230] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 162 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 162, 'op': 'addl'}
    instructions[4231] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 162 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 162, 'op': 'load'}
    instructions[4232] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 162 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 162, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4233] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 162 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 162, 'op': 'load'}
    instructions[4234] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 162 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 162, 'op': 'add'}
    instructions[4235] = {5'd1, 4'd2, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 162 {'a': 4, 'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 162, 'op': 'addl'}
    instructions[4236] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 162 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 162, 'op': 'store'}
    instructions[4237] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164, 'op': 'literal'}
    instructions[4238] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164, 'op': 'store'}
    instructions[4239] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164, 'op': 'addl'}
    instructions[4240] = {5'd1, 4'd8, 4'd4, 16'd1465};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164 {'a': 4, 'literal': 1465, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164, 'op': 'addl'}
    instructions[4241] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164, 'op': 'addl'}
    instructions[4242] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164, 'op': 'load'}
    instructions[4243] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4244] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164, 'op': 'load'}
    instructions[4245] = {5'd10, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164, 'op': 'and'}
    instructions[4246] = {5'd8, 4'd0, 4'd8, 16'd4264};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164 {'a': 8, 'label': 4264, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164, 'op': 'jmp_if_false'}
    instructions[4247] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164, 'op': 'literal'}
    instructions[4248] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164, 'op': 'store'}
    instructions[4249] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164, 'op': 'addl'}
    instructions[4250] = {5'd1, 4'd8, 4'd4, 16'd1469};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164 {'a': 4, 'literal': 1469, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164, 'op': 'addl'}
    instructions[4251] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164, 'op': 'store'}
    instructions[4252] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164, 'op': 'addl'}
    instructions[4253] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164, 'op': 'addl'}
    instructions[4254] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164, 'op': 'addl'}
    instructions[4255] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164, 'op': 'load'}
    instructions[4256] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4257] = {5'd5, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164, 'op': 'load'}
    instructions[4258] = {5'd11, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164, 'op': 'add'}
    instructions[4259] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164, 'op': 'addl'}
    instructions[4260] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4261] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164, 'op': 'load'}
    instructions[4262] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164, 'op': 'store'}
    instructions[4263] = {5'd12, 4'd0, 4'd0, 16'd4280};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164 {'label': 4280, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 164, 'op': 'goto'}
    instructions[4264] = {5'd0, 4'd8, 4'd0, 16'd49};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 165 {'literal': 49, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 165, 'op': 'literal'}
    instructions[4265] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 165 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 165, 'op': 'store'}
    instructions[4266] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 165 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 165, 'op': 'addl'}
    instructions[4267] = {5'd1, 4'd8, 4'd4, 16'd1469};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 165 {'a': 4, 'literal': 1469, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 165, 'op': 'addl'}
    instructions[4268] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 165 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 165, 'op': 'store'}
    instructions[4269] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 165 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 165, 'op': 'addl'}
    instructions[4270] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 165 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 165, 'op': 'addl'}
    instructions[4271] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 165 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 165, 'op': 'addl'}
    instructions[4272] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 165 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 165, 'op': 'load'}
    instructions[4273] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 165 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 165, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4274] = {5'd5, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 165 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 165, 'op': 'load'}
    instructions[4275] = {5'd11, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 165 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 165, 'op': 'add'}
    instructions[4276] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 165 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 165, 'op': 'addl'}
    instructions[4277] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 165 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 165, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4278] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 165 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 165, 'op': 'load'}
    instructions[4279] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 165 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 165, 'op': 'store'}
    instructions[4280] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 166 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 166, 'op': 'addl'}
    instructions[4281] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 166 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 166, 'op': 'addl'}
    instructions[4282] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 166 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 166, 'op': 'load'}
    instructions[4283] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 166 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 166, 'op': 'store'}
    instructions[4284] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 166 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 166, 'op': 'addl'}
    instructions[4285] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 166 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 166, 'op': 'literal'}
    instructions[4286] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 166 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 166, 'op': 'store'}
    instructions[4287] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 166 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 166, 'op': 'addl'}
    instructions[4288] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 166 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 166, 'op': 'addl'}
    instructions[4289] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 166 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 166, 'op': 'addl'}
    instructions[4290] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 166 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 166, 'op': 'load'}
    instructions[4291] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 166 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 166, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4292] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 166 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 166, 'op': 'load'}
    instructions[4293] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 166 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 166, 'op': 'add'}
    instructions[4294] = {5'd1, 4'd2, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 166 {'a': 4, 'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 166, 'op': 'addl'}
    instructions[4295] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 166 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 166, 'op': 'store'}
    instructions[4296] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 166 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 166, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4297] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 166 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 166, 'op': 'load'}
    instructions[4298] = {5'd0, 4'd8, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167 {'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167, 'op': 'literal'}
    instructions[4299] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167, 'op': 'store'}
    instructions[4300] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167, 'op': 'addl'}
    instructions[4301] = {5'd1, 4'd8, 4'd4, 16'd1465};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167 {'a': 4, 'literal': 1465, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167, 'op': 'addl'}
    instructions[4302] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167, 'op': 'addl'}
    instructions[4303] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167, 'op': 'load'}
    instructions[4304] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4305] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167, 'op': 'load'}
    instructions[4306] = {5'd10, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167, 'op': 'and'}
    instructions[4307] = {5'd8, 4'd0, 4'd8, 16'd4325};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167 {'a': 8, 'label': 4325, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167, 'op': 'jmp_if_false'}
    instructions[4308] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167, 'op': 'literal'}
    instructions[4309] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167, 'op': 'store'}
    instructions[4310] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167, 'op': 'addl'}
    instructions[4311] = {5'd1, 4'd8, 4'd4, 16'd1469};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167 {'a': 4, 'literal': 1469, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167, 'op': 'addl'}
    instructions[4312] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167, 'op': 'store'}
    instructions[4313] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167, 'op': 'addl'}
    instructions[4314] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167, 'op': 'addl'}
    instructions[4315] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167, 'op': 'addl'}
    instructions[4316] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167, 'op': 'load'}
    instructions[4317] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4318] = {5'd5, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167, 'op': 'load'}
    instructions[4319] = {5'd11, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167, 'op': 'add'}
    instructions[4320] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167, 'op': 'addl'}
    instructions[4321] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4322] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167, 'op': 'load'}
    instructions[4323] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167, 'op': 'store'}
    instructions[4324] = {5'd12, 4'd0, 4'd0, 16'd4341};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167 {'label': 4341, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 167, 'op': 'goto'}
    instructions[4325] = {5'd0, 4'd8, 4'd0, 16'd49};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 168 {'literal': 49, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 168, 'op': 'literal'}
    instructions[4326] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 168 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 168, 'op': 'store'}
    instructions[4327] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 168 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 168, 'op': 'addl'}
    instructions[4328] = {5'd1, 4'd8, 4'd4, 16'd1469};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 168 {'a': 4, 'literal': 1469, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 168, 'op': 'addl'}
    instructions[4329] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 168 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 168, 'op': 'store'}
    instructions[4330] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 168 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 168, 'op': 'addl'}
    instructions[4331] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 168 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 168, 'op': 'addl'}
    instructions[4332] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 168 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 168, 'op': 'addl'}
    instructions[4333] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 168 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 168, 'op': 'load'}
    instructions[4334] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 168 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 168, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4335] = {5'd5, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 168 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 168, 'op': 'load'}
    instructions[4336] = {5'd11, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 168 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 168, 'op': 'add'}
    instructions[4337] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 168 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 168, 'op': 'addl'}
    instructions[4338] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 168 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 168, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4339] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 168 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 168, 'op': 'load'}
    instructions[4340] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 168 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 168, 'op': 'store'}
    instructions[4341] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 169 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 169, 'op': 'addl'}
    instructions[4342] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 169 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 169, 'op': 'addl'}
    instructions[4343] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 169 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 169, 'op': 'load'}
    instructions[4344] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 169 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 169, 'op': 'store'}
    instructions[4345] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 169 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 169, 'op': 'addl'}
    instructions[4346] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 169 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 169, 'op': 'literal'}
    instructions[4347] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 169 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 169, 'op': 'store'}
    instructions[4348] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 169 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 169, 'op': 'addl'}
    instructions[4349] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 169 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 169, 'op': 'addl'}
    instructions[4350] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 169 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 169, 'op': 'addl'}
    instructions[4351] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 169 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 169, 'op': 'load'}
    instructions[4352] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 169 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 169, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4353] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 169 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 169, 'op': 'load'}
    instructions[4354] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 169 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 169, 'op': 'add'}
    instructions[4355] = {5'd1, 4'd2, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 169 {'a': 4, 'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 169, 'op': 'addl'}
    instructions[4356] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 169 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 169, 'op': 'store'}
    instructions[4357] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 169 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 169, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4358] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 169 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 169, 'op': 'load'}
    instructions[4359] = {5'd0, 4'd8, 4'd0, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170 {'literal': 4, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170, 'op': 'literal'}
    instructions[4360] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170, 'op': 'store'}
    instructions[4361] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170, 'op': 'addl'}
    instructions[4362] = {5'd1, 4'd8, 4'd4, 16'd1465};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170 {'a': 4, 'literal': 1465, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170, 'op': 'addl'}
    instructions[4363] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170, 'op': 'addl'}
    instructions[4364] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170, 'op': 'load'}
    instructions[4365] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4366] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170, 'op': 'load'}
    instructions[4367] = {5'd10, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170, 'op': 'and'}
    instructions[4368] = {5'd8, 4'd0, 4'd8, 16'd4386};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170 {'a': 8, 'label': 4386, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170, 'op': 'jmp_if_false'}
    instructions[4369] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170, 'op': 'literal'}
    instructions[4370] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170, 'op': 'store'}
    instructions[4371] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170, 'op': 'addl'}
    instructions[4372] = {5'd1, 4'd8, 4'd4, 16'd1469};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170 {'a': 4, 'literal': 1469, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170, 'op': 'addl'}
    instructions[4373] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170, 'op': 'store'}
    instructions[4374] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170, 'op': 'addl'}
    instructions[4375] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170, 'op': 'addl'}
    instructions[4376] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170, 'op': 'addl'}
    instructions[4377] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170, 'op': 'load'}
    instructions[4378] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4379] = {5'd5, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170, 'op': 'load'}
    instructions[4380] = {5'd11, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170, 'op': 'add'}
    instructions[4381] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170, 'op': 'addl'}
    instructions[4382] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4383] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170, 'op': 'load'}
    instructions[4384] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170, 'op': 'store'}
    instructions[4385] = {5'd12, 4'd0, 4'd0, 16'd4402};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170 {'label': 4402, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 170, 'op': 'goto'}
    instructions[4386] = {5'd0, 4'd8, 4'd0, 16'd49};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 171 {'literal': 49, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 171, 'op': 'literal'}
    instructions[4387] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 171 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 171, 'op': 'store'}
    instructions[4388] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 171 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 171, 'op': 'addl'}
    instructions[4389] = {5'd1, 4'd8, 4'd4, 16'd1469};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 171 {'a': 4, 'literal': 1469, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 171, 'op': 'addl'}
    instructions[4390] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 171 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 171, 'op': 'store'}
    instructions[4391] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 171 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 171, 'op': 'addl'}
    instructions[4392] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 171 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 171, 'op': 'addl'}
    instructions[4393] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 171 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 171, 'op': 'addl'}
    instructions[4394] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 171 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 171, 'op': 'load'}
    instructions[4395] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 171 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 171, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4396] = {5'd5, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 171 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 171, 'op': 'load'}
    instructions[4397] = {5'd11, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 171 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 171, 'op': 'add'}
    instructions[4398] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 171 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 171, 'op': 'addl'}
    instructions[4399] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 171 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 171, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4400] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 171 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 171, 'op': 'load'}
    instructions[4401] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 171 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 171, 'op': 'store'}
    instructions[4402] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 172 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 172, 'op': 'addl'}
    instructions[4403] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 172 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 172, 'op': 'addl'}
    instructions[4404] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 172 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 172, 'op': 'load'}
    instructions[4405] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 172 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 172, 'op': 'store'}
    instructions[4406] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 172 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 172, 'op': 'addl'}
    instructions[4407] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 172 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 172, 'op': 'literal'}
    instructions[4408] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 172 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 172, 'op': 'store'}
    instructions[4409] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 172 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 172, 'op': 'addl'}
    instructions[4410] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 172 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 172, 'op': 'addl'}
    instructions[4411] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 172 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 172, 'op': 'addl'}
    instructions[4412] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 172 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 172, 'op': 'load'}
    instructions[4413] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 172 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 172, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4414] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 172 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 172, 'op': 'load'}
    instructions[4415] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 172 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 172, 'op': 'add'}
    instructions[4416] = {5'd1, 4'd2, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 172 {'a': 4, 'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 172, 'op': 'addl'}
    instructions[4417] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 172 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 172, 'op': 'store'}
    instructions[4418] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 172 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 172, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4419] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 172 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 172, 'op': 'load'}
    instructions[4420] = {5'd0, 4'd8, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173 {'literal': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173, 'op': 'literal'}
    instructions[4421] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173, 'op': 'store'}
    instructions[4422] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173, 'op': 'addl'}
    instructions[4423] = {5'd1, 4'd8, 4'd4, 16'd1465};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173 {'a': 4, 'literal': 1465, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173, 'op': 'addl'}
    instructions[4424] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173, 'op': 'addl'}
    instructions[4425] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173, 'op': 'load'}
    instructions[4426] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4427] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173, 'op': 'load'}
    instructions[4428] = {5'd10, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173, 'op': 'and'}
    instructions[4429] = {5'd8, 4'd0, 4'd8, 16'd4447};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173 {'a': 8, 'label': 4447, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173, 'op': 'jmp_if_false'}
    instructions[4430] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173, 'op': 'literal'}
    instructions[4431] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173, 'op': 'store'}
    instructions[4432] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173, 'op': 'addl'}
    instructions[4433] = {5'd1, 4'd8, 4'd4, 16'd1469};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173 {'a': 4, 'literal': 1469, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173, 'op': 'addl'}
    instructions[4434] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173, 'op': 'store'}
    instructions[4435] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173, 'op': 'addl'}
    instructions[4436] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173, 'op': 'addl'}
    instructions[4437] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173, 'op': 'addl'}
    instructions[4438] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173, 'op': 'load'}
    instructions[4439] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4440] = {5'd5, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173, 'op': 'load'}
    instructions[4441] = {5'd11, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173, 'op': 'add'}
    instructions[4442] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173, 'op': 'addl'}
    instructions[4443] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4444] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173, 'op': 'load'}
    instructions[4445] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173, 'op': 'store'}
    instructions[4446] = {5'd12, 4'd0, 4'd0, 16'd4463};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173 {'label': 4463, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 173, 'op': 'goto'}
    instructions[4447] = {5'd0, 4'd8, 4'd0, 16'd49};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 174 {'literal': 49, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 174, 'op': 'literal'}
    instructions[4448] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 174 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 174, 'op': 'store'}
    instructions[4449] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 174 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 174, 'op': 'addl'}
    instructions[4450] = {5'd1, 4'd8, 4'd4, 16'd1469};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 174 {'a': 4, 'literal': 1469, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 174, 'op': 'addl'}
    instructions[4451] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 174 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 174, 'op': 'store'}
    instructions[4452] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 174 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 174, 'op': 'addl'}
    instructions[4453] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 174 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 174, 'op': 'addl'}
    instructions[4454] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 174 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 174, 'op': 'addl'}
    instructions[4455] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 174 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 174, 'op': 'load'}
    instructions[4456] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 174 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 174, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4457] = {5'd5, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 174 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 174, 'op': 'load'}
    instructions[4458] = {5'd11, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 174 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 174, 'op': 'add'}
    instructions[4459] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 174 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 174, 'op': 'addl'}
    instructions[4460] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 174 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 174, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4461] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 174 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 174, 'op': 'load'}
    instructions[4462] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 174 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 174, 'op': 'store'}
    instructions[4463] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 176 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 176, 'op': 'store'}
    instructions[4464] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 176 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 176, 'op': 'addl'}
    instructions[4465] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 176 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 176, 'op': 'store'}
    instructions[4466] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 176 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 176, 'op': 'addl'}
    instructions[4467] = {5'd1, 4'd8, 4'd4, 16'd1469};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 176 {'a': 4, 'literal': 1469, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 176, 'op': 'addl'}
    instructions[4468] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 176 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 176, 'op': 'store'}
    instructions[4469] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 176 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 176, 'op': 'addl'}
    instructions[4470] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 176 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 176, 'op': 'addl'}
    instructions[4471] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 176 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 176, 'op': 'addl'}
    instructions[4472] = {5'd3, 4'd6, 4'd0, 16'd4685};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 176 {'z': 6, 'label': 4685, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 176, 'op': 'call'}
    instructions[4473] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 176 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 176, 'op': 'addl'}
    instructions[4474] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 176 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 176, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4475] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 176 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 176, 'op': 'load'}
    instructions[4476] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 176 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 176, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4477] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 176 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 176, 'op': 'load'}
    instructions[4478] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 176 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 176, 'op': 'addl'}
    instructions[4479] = {5'd12, 4'd0, 4'd0, 16'd4493};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 107 {'label': 4493, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 107, 'op': 'goto'}
    instructions[4480] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 178 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 178, 'op': 'store'}
    instructions[4481] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 178 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 178, 'op': 'addl'}
    instructions[4482] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 178 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 178, 'op': 'store'}
    instructions[4483] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 178 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 178, 'op': 'addl'}
    instructions[4484] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 178 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 178, 'op': 'addl'}
    instructions[4485] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 178 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 178, 'op': 'addl'}
    instructions[4486] = {5'd3, 4'd6, 4'd0, 16'd6172};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 178 {'z': 6, 'label': 6172, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 178, 'op': 'call'}
    instructions[4487] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 178 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 178, 'op': 'addl'}
    instructions[4488] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 178 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 178, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4489] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 178 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 178, 'op': 'load'}
    instructions[4490] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 178 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 178, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4491] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 178 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 178, 'op': 'load'}
    instructions[4492] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 178 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 178, 'op': 'addl'}
    instructions[4493] = {5'd12, 4'd0, 4'd0, 16'd2981};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 92 {'label': 2981, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 92, 'op': 'goto'}
    instructions[4494] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 49 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 49, 'op': 'addl'}
    instructions[4495] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 49 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 49, 'op': 'addl'}
    instructions[4496] = {5'd19, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 49 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 49, 'op': 'return'}
    instructions[4497] = {5'd1, 4'd3, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73 {'a': 3, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73, 'op': 'addl'}
    instructions[4498] = {5'd2, 4'd0, 4'd3, 16'd6};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'store'}
    instructions[4499] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[4500] = {5'd2, 4'd0, 4'd3, 16'd7};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'store'}
    instructions[4501] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[4502] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[4503] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[4504] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'load'}
    instructions[4505] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'store'}
    instructions[4506] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[4507] = {5'd0, 4'd8, 4'd0, 16'd7};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'literal': 7, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'literal'}
    instructions[4508] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[4509] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'load'}
    instructions[4510] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'store'}
    instructions[4511] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[4512] = {5'd1, 4'd7, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 4, 'literal': 0, 'z': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[4513] = {5'd1, 4'd4, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[4514] = {5'd3, 4'd6, 4'd0, 16'd4524};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'z': 6, 'label': 4524, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'call'}
    instructions[4515] = {5'd1, 4'd3, 4'd3, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': -2, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[4516] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4517] = {5'd5, 4'd7, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'z': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'load'}
    instructions[4518] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4519] = {5'd5, 4'd6, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'z': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'load'}
    instructions[4520] = {5'd1, 4'd3, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[4521] = {5'd1, 4'd3, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73 {'a': 4, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73, 'op': 'addl'}
    instructions[4522] = {5'd1, 4'd4, 4'd7, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73 {'a': 7, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73, 'op': 'addl'}
    instructions[4523] = {5'd19, 4'd0, 4'd6, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73 {'a': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73, 'op': 'return'}
    instructions[4524] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23, 'op': 'addl'}
    instructions[4525] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 24 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 24, 'op': 'literal'}
    instructions[4526] = {5'd1, 4'd2, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 24 {'a': 4, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 24, 'op': 'addl'}
    instructions[4527] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 24 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 24, 'op': 'store'}
    instructions[4528] = {5'd1, 4'd8, 4'd4, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 4, 'literal': -2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'addl'}
    instructions[4529] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'addl'}
    instructions[4530] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'load'}
    instructions[4531] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'store'}
    instructions[4532] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'addl'}
    instructions[4533] = {5'd1, 4'd8, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 4, 'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'addl'}
    instructions[4534] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'addl'}
    instructions[4535] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'load'}
    instructions[4536] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4537] = {5'd5, 4'd2, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 3, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'load'}
    instructions[4538] = {5'd11, 4'd8, 4'd8, 16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 8, 'z': 8, 'b': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'add'}
    instructions[4539] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'addl'}
    instructions[4540] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'load'}
    instructions[4541] = {5'd8, 4'd0, 4'd8, 16'd4583};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 29 {'a': 8, 'label': 4583, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 29, 'op': 'jmp_if_false'}
    instructions[4542] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[4543] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[4544] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'load'}
    instructions[4545] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'store'}
    instructions[4546] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[4547] = {5'd1, 4'd8, 4'd4, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 4, 'literal': -2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[4548] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[4549] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'load'}
    instructions[4550] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'store'}
    instructions[4551] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[4552] = {5'd1, 4'd8, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 4, 'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[4553] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[4554] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'load'}
    instructions[4555] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4556] = {5'd5, 4'd2, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'load'}
    instructions[4557] = {5'd11, 4'd8, 4'd8, 16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 8, 'z': 8, 'b': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'add'}
    instructions[4558] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[4559] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'load'}
    instructions[4560] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4561] = {5'd5, 4'd0, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'z': 0, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'load'}
    instructions[4562] = {5'd17, 4'd0, 4'd0, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 0, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'write'}
    instructions[4563] = {5'd1, 4'd3, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[4564] = {5'd1, 4'd8, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 4, 'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[4565] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[4566] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'load'}
    instructions[4567] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'store'}
    instructions[4568] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[4569] = {5'd0, 4'd8, 4'd0, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'literal': 1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'literal'}
    instructions[4570] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'store'}
    instructions[4571] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[4572] = {5'd1, 4'd8, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 4, 'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[4573] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[4574] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'load'}
    instructions[4575] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4576] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'load'}
    instructions[4577] = {5'd11, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'add'}
    instructions[4578] = {5'd1, 4'd2, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 4, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[4579] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'store'}
    instructions[4580] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4581] = {5'd5, 4'd8, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'load'}
    instructions[4582] = {5'd12, 4'd0, 4'd0, 16'd4584};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 29 {'label': 4584, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 29, 'op': 'goto'}
    instructions[4583] = {5'd12, 4'd0, 4'd0, 16'd4585};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 29 {'label': 4585, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 29, 'op': 'goto'}
    instructions[4584] = {5'd12, 4'd0, 4'd0, 16'd4528};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'label': 4528, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'goto'}
    instructions[4585] = {5'd1, 4'd3, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23 {'a': 4, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23, 'op': 'addl'}
    instructions[4586] = {5'd1, 4'd4, 4'd7, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23 {'a': 7, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23, 'op': 'addl'}
    instructions[4587] = {5'd19, 4'd0, 4'd6, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23 {'a': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23, 'op': 'return'}
    instructions[4588] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 39 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 39, 'op': 'addl'}
    instructions[4589] = {5'd1, 4'd8, 4'd4, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 40 {'a': 4, 'literal': -2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 40, 'op': 'addl'}
    instructions[4590] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 40 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 40, 'op': 'addl'}
    instructions[4591] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 40 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 40, 'op': 'load'}
    instructions[4592] = {5'd1, 4'd2, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 40 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 40, 'op': 'addl'}
    instructions[4593] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 40 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 40, 'op': 'store'}
    instructions[4594] = {5'd1, 4'd8, 4'd4, -16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 41 {'a': 4, 'literal': -4, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 41, 'op': 'addl'}
    instructions[4595] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 41 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 41, 'op': 'addl'}
    instructions[4596] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 41 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 41, 'op': 'load'}
    instructions[4597] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 41 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 41, 'op': 'store'}
    instructions[4598] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 41 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 41, 'op': 'addl'}
    instructions[4599] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 41 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 41, 'op': 'addl'}
    instructions[4600] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 41 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 41, 'op': 'addl'}
    instructions[4601] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 41 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 41, 'op': 'load'}
    instructions[4602] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 41 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 41, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4603] = {5'd5, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 41 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 41, 'op': 'load'}
    instructions[4604] = {5'd11, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 41 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 41, 'op': 'add'}
    instructions[4605] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 41 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 41, 'op': 'addl'}
    instructions[4606] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 41 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 41, 'op': 'load'}
    instructions[4607] = {5'd8, 4'd0, 4'd8, 16'd4677};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 46 {'a': 8, 'label': 4677, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 46, 'op': 'jmp_if_false'}
    instructions[4608] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 42 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 42, 'op': 'addl'}
    instructions[4609] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 42 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 42, 'op': 'addl'}
    instructions[4610] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 42 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 42, 'op': 'load'}
    instructions[4611] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 42 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 42, 'op': 'store'}
    instructions[4612] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 42 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 42, 'op': 'addl'}
    instructions[4613] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 42 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 42, 'op': 'addl'}
    instructions[4614] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 42 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 42, 'op': 'addl'}
    instructions[4615] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 42 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 42, 'op': 'load'}
    instructions[4616] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 42 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 42, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4617] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 42 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 42, 'op': 'load'}
    instructions[4618] = {5'd13, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 42 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 42, 'op': 'equal'}
    instructions[4619] = {5'd8, 4'd0, 4'd8, 16'd4627};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 42 {'a': 8, 'label': 4627, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 42, 'op': 'jmp_if_false'}
    instructions[4620] = {5'd0, 4'd8, 4'd0, 16'd65535};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 42 {'literal': 65535, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 42, 'op': 'literal'}
    instructions[4621] = {5'd0, 4'd2, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 42 {'literal': 6, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 42, 'op': 'literal'}
    instructions[4622] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 42 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 42, 'op': 'store'}
    instructions[4623] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 42 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 42, 'op': 'addl'}
    instructions[4624] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 42 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 42, 'op': 'addl'}
    instructions[4625] = {5'd19, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 42 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 42, 'op': 'return'}
    instructions[4626] = {5'd12, 4'd0, 4'd0, 16'd4627};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 42 {'label': 4627, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 42, 'op': 'goto'}
    instructions[4627] = {5'd1, 4'd8, 4'd4, -16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43 {'a': 4, 'literal': -3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43, 'op': 'addl'}
    instructions[4628] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43, 'op': 'addl'}
    instructions[4629] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43, 'op': 'load'}
    instructions[4630] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43, 'op': 'store'}
    instructions[4631] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43, 'op': 'addl'}
    instructions[4632] = {5'd1, 4'd8, 4'd4, -16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43 {'a': 4, 'literal': -4, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43, 'op': 'addl'}
    instructions[4633] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43, 'op': 'addl'}
    instructions[4634] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43, 'op': 'load'}
    instructions[4635] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43, 'op': 'store'}
    instructions[4636] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43, 'op': 'addl'}
    instructions[4637] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43, 'op': 'addl'}
    instructions[4638] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43, 'op': 'addl'}
    instructions[4639] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43, 'op': 'load'}
    instructions[4640] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4641] = {5'd5, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43, 'op': 'load'}
    instructions[4642] = {5'd11, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43, 'op': 'add'}
    instructions[4643] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43, 'op': 'addl'}
    instructions[4644] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43, 'op': 'load'}
    instructions[4645] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4646] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43, 'op': 'load'}
    instructions[4647] = {5'd13, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43, 'op': 'equal'}
    instructions[4648] = {5'd8, 4'd0, 4'd8, 16'd4658};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43 {'a': 8, 'label': 4658, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43, 'op': 'jmp_if_false'}
    instructions[4649] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43, 'op': 'addl'}
    instructions[4650] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43, 'op': 'addl'}
    instructions[4651] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43, 'op': 'load'}
    instructions[4652] = {5'd0, 4'd2, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43 {'literal': 6, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43, 'op': 'literal'}
    instructions[4653] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43, 'op': 'store'}
    instructions[4654] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43, 'op': 'addl'}
    instructions[4655] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43, 'op': 'addl'}
    instructions[4656] = {5'd19, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43, 'op': 'return'}
    instructions[4657] = {5'd12, 4'd0, 4'd0, 16'd4658};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43 {'label': 4658, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 43, 'op': 'goto'}
    instructions[4658] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 44 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 44, 'op': 'addl'}
    instructions[4659] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 44 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 44, 'op': 'addl'}
    instructions[4660] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 44 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 44, 'op': 'load'}
    instructions[4661] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 44 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 44, 'op': 'store'}
    instructions[4662] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 44 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 44, 'op': 'addl'}
    instructions[4663] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 44 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 44, 'op': 'literal'}
    instructions[4664] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 44 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 44, 'op': 'store'}
    instructions[4665] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 44 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 44, 'op': 'addl'}
    instructions[4666] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 44 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 44, 'op': 'addl'}
    instructions[4667] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 44 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 44, 'op': 'addl'}
    instructions[4668] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 44 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 44, 'op': 'load'}
    instructions[4669] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 44 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 44, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4670] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 44 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 44, 'op': 'load'}
    instructions[4671] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 44 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 44, 'op': 'add'}
    instructions[4672] = {5'd1, 4'd2, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 44 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 44, 'op': 'addl'}
    instructions[4673] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 44 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 44, 'op': 'store'}
    instructions[4674] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 44 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 44, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4675] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 44 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 44, 'op': 'load'}
    instructions[4676] = {5'd12, 4'd0, 4'd0, 16'd4678};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 46 {'label': 4678, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 46, 'op': 'goto'}
    instructions[4677] = {5'd12, 4'd0, 4'd0, 16'd4679};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 46 {'label': 4679, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 46, 'op': 'goto'}
    instructions[4678] = {5'd12, 4'd0, 4'd0, 16'd4594};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 41 {'label': 4594, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 41, 'op': 'goto'}
    instructions[4679] = {5'd0, 4'd8, 4'd0, 16'd65535};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 46 {'literal': 65535, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 46, 'op': 'literal'}
    instructions[4680] = {5'd0, 4'd2, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 46 {'literal': 6, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 46, 'op': 'literal'}
    instructions[4681] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 46 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 46, 'op': 'store'}
    instructions[4682] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 46 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 46, 'op': 'addl'}
    instructions[4683] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 46 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 46, 'op': 'addl'}
    instructions[4684] = {5'd19, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 46 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 46, 'op': 'return'}
    instructions[4685] = {5'd1, 4'd3, 4'd3, 16'd124};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 106 {'a': 3, 'literal': 124, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 106, 'op': 'addl'}
    instructions[4686] = {5'd0, 4'd8, 4'd0, 16'd72};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 72, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4687] = {5'd1, 4'd2, 4'd4, 16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 5, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4688] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4689] = {5'd0, 4'd8, 4'd0, 16'd84};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 84, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4690] = {5'd1, 4'd2, 4'd4, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 6, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4691] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4692] = {5'd0, 4'd8, 4'd0, 16'd84};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 84, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4693] = {5'd1, 4'd2, 4'd4, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 7, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4694] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4695] = {5'd0, 4'd8, 4'd0, 16'd80};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 80, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4696] = {5'd1, 4'd2, 4'd4, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 8, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4697] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4698] = {5'd0, 4'd8, 4'd0, 16'd47};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 47, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4699] = {5'd1, 4'd2, 4'd4, 16'd9};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 9, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4700] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4701] = {5'd0, 4'd8, 4'd0, 16'd49};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 49, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4702] = {5'd1, 4'd2, 4'd4, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 10, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4703] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4704] = {5'd0, 4'd8, 4'd0, 16'd46};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 46, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4705] = {5'd1, 4'd2, 4'd4, 16'd11};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 11, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4706] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4707] = {5'd0, 4'd8, 4'd0, 16'd49};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 49, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4708] = {5'd1, 4'd2, 4'd4, 16'd12};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 12, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4709] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4710] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4711] = {5'd1, 4'd2, 4'd4, 16'd13};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 13, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4712] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4713] = {5'd0, 4'd8, 4'd0, 16'd50};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 50, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4714] = {5'd1, 4'd2, 4'd4, 16'd14};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 14, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4715] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4716] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4717] = {5'd1, 4'd2, 4'd4, 16'd15};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 15, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4718] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4719] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4720] = {5'd1, 4'd2, 4'd4, 16'd16};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 16, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4721] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4722] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4723] = {5'd1, 4'd2, 4'd4, 16'd17};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 17, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4724] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4725] = {5'd0, 4'd8, 4'd0, 16'd79};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 79, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4726] = {5'd1, 4'd2, 4'd4, 16'd18};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 18, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4727] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4728] = {5'd0, 4'd8, 4'd0, 16'd75};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 75, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4729] = {5'd1, 4'd2, 4'd4, 16'd19};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 19, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4730] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4731] = {5'd0, 4'd8, 4'd0, 16'd13};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 13, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4732] = {5'd1, 4'd2, 4'd4, 16'd20};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 20, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4733] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4734] = {5'd0, 4'd8, 4'd0, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 10, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4735] = {5'd1, 4'd2, 4'd4, 16'd21};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 21, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4736] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4737] = {5'd0, 4'd8, 4'd0, 16'd68};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 68, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4738] = {5'd1, 4'd2, 4'd4, 16'd22};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 22, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4739] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4740] = {5'd0, 4'd8, 4'd0, 16'd97};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 97, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4741] = {5'd1, 4'd2, 4'd4, 16'd23};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 23, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4742] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4743] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4744] = {5'd1, 4'd2, 4'd4, 16'd24};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 24, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4745] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4746] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4747] = {5'd1, 4'd2, 4'd4, 16'd25};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 25, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4748] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4749] = {5'd0, 4'd8, 4'd0, 16'd58};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 58, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4750] = {5'd1, 4'd2, 4'd4, 16'd26};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 26, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4751] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4752] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4753] = {5'd1, 4'd2, 4'd4, 16'd27};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 27, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4754] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4755] = {5'd0, 4'd8, 4'd0, 16'd84};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 84, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4756] = {5'd1, 4'd2, 4'd4, 16'd28};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 28, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4757] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4758] = {5'd0, 4'd8, 4'd0, 16'd104};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 104, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4759] = {5'd1, 4'd2, 4'd4, 16'd29};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 29, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4760] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4761] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4762] = {5'd1, 4'd2, 4'd4, 16'd30};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 30, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4763] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4764] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4765] = {5'd1, 4'd2, 4'd4, 16'd31};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 31, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4766] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4767] = {5'd0, 4'd8, 4'd0, 16'd79};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 79, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4768] = {5'd1, 4'd2, 4'd4, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 32, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4769] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4770] = {5'd0, 4'd8, 4'd0, 16'd99};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 99, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4771] = {5'd1, 4'd2, 4'd4, 16'd33};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 33, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4772] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4773] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4774] = {5'd1, 4'd2, 4'd4, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 34, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4775] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4776] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4777] = {5'd1, 4'd2, 4'd4, 16'd35};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 35, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4778] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4779] = {5'd0, 4'd8, 4'd0, 16'd51};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 51, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4780] = {5'd1, 4'd2, 4'd4, 16'd36};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 36, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4781] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4782] = {5'd0, 4'd8, 4'd0, 16'd49};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 49, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4783] = {5'd1, 4'd2, 4'd4, 16'd37};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 37, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4784] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4785] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4786] = {5'd1, 4'd2, 4'd4, 16'd38};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 38, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4787] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4788] = {5'd0, 4'd8, 4'd0, 16'd49};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 49, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4789] = {5'd1, 4'd2, 4'd4, 16'd39};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 39, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4790] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4791] = {5'd0, 4'd8, 4'd0, 16'd57};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 57, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4792] = {5'd1, 4'd2, 4'd4, 16'd40};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 40, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4793] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4794] = {5'd0, 4'd8, 4'd0, 16'd58};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 58, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4795] = {5'd1, 4'd2, 4'd4, 16'd41};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 41, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4796] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4797] = {5'd0, 4'd8, 4'd0, 16'd49};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 49, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4798] = {5'd1, 4'd2, 4'd4, 16'd42};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 42, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4799] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4800] = {5'd0, 4'd8, 4'd0, 16'd54};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 54, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4801] = {5'd1, 4'd2, 4'd4, 16'd43};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 43, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4802] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4803] = {5'd0, 4'd8, 4'd0, 16'd58};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 58, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4804] = {5'd1, 4'd2, 4'd4, 16'd44};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 44, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4805] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4806] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4807] = {5'd1, 4'd2, 4'd4, 16'd45};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 45, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4808] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4809] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4810] = {5'd1, 4'd2, 4'd4, 16'd46};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 46, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4811] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4812] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4813] = {5'd1, 4'd2, 4'd4, 16'd47};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 47, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4814] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4815] = {5'd0, 4'd8, 4'd0, 16'd50};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 50, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4816] = {5'd1, 4'd2, 4'd4, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 48, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4817] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4818] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4819] = {5'd1, 4'd2, 4'd4, 16'd49};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 49, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4820] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4821] = {5'd0, 4'd8, 4'd0, 16'd49};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 49, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4822] = {5'd1, 4'd2, 4'd4, 16'd50};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 50, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4823] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4824] = {5'd0, 4'd8, 4'd0, 16'd51};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 51, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4825] = {5'd1, 4'd2, 4'd4, 16'd51};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 51, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4826] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4827] = {5'd0, 4'd8, 4'd0, 16'd13};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 13, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4828] = {5'd1, 4'd2, 4'd4, 16'd52};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 52, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4829] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4830] = {5'd0, 4'd8, 4'd0, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 10, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4831] = {5'd1, 4'd2, 4'd4, 16'd53};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 53, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4832] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4833] = {5'd0, 4'd8, 4'd0, 16'd83};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 83, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4834] = {5'd1, 4'd2, 4'd4, 16'd54};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 54, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4835] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4836] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4837] = {5'd1, 4'd2, 4'd4, 16'd55};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 55, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4838] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4839] = {5'd0, 4'd8, 4'd0, 16'd114};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 114, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4840] = {5'd1, 4'd2, 4'd4, 16'd56};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 56, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4841] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4842] = {5'd0, 4'd8, 4'd0, 16'd118};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 118, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4843] = {5'd1, 4'd2, 4'd4, 16'd57};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 57, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4844] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4845] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4846] = {5'd1, 4'd2, 4'd4, 16'd58};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 58, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4847] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4848] = {5'd0, 4'd8, 4'd0, 16'd114};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 114, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4849] = {5'd1, 4'd2, 4'd4, 16'd59};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 59, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4850] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4851] = {5'd0, 4'd8, 4'd0, 16'd58};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 58, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4852] = {5'd1, 4'd2, 4'd4, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 60, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4853] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4854] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4855] = {5'd1, 4'd2, 4'd4, 16'd61};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 61, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4856] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4857] = {5'd0, 4'd8, 4'd0, 16'd99};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 99, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4858] = {5'd1, 4'd2, 4'd4, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 62, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4859] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4860] = {5'd0, 4'd8, 4'd0, 16'd104};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 104, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4861] = {5'd1, 4'd2, 4'd4, 16'd63};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 63, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4862] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4863] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4864] = {5'd1, 4'd2, 4'd4, 16'd64};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 64, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4865] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4866] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4867] = {5'd1, 4'd2, 4'd4, 16'd65};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 65, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4868] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4869] = {5'd0, 4'd8, 4'd0, 16'd115};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 115, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4870] = {5'd1, 4'd2, 4'd4, 16'd66};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 66, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4871] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4872] = {5'd0, 4'd8, 4'd0, 16'd45};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 45, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4873] = {5'd1, 4'd2, 4'd4, 16'd67};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 67, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4874] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4875] = {5'd0, 4'd8, 4'd0, 16'd119};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 119, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4876] = {5'd1, 4'd2, 4'd4, 16'd68};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 68, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4877] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4878] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4879] = {5'd1, 4'd2, 4'd4, 16'd69};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 69, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4880] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4881] = {5'd0, 4'd8, 4'd0, 16'd98};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 98, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4882] = {5'd1, 4'd2, 4'd4, 16'd70};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 70, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4883] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4884] = {5'd0, 4'd8, 4'd0, 16'd47};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 47, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4885] = {5'd1, 4'd2, 4'd4, 16'd71};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 71, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4886] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4887] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4888] = {5'd1, 4'd2, 4'd4, 16'd72};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 72, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4889] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4890] = {5'd0, 4'd8, 4'd0, 16'd46};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 46, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4891] = {5'd1, 4'd2, 4'd4, 16'd73};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 73, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4892] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4893] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4894] = {5'd1, 4'd2, 4'd4, 16'd74};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 74, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4895] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4896] = {5'd0, 4'd8, 4'd0, 16'd13};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 13, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4897] = {5'd1, 4'd2, 4'd4, 16'd75};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 75, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4898] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4899] = {5'd0, 4'd8, 4'd0, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 10, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4900] = {5'd1, 4'd2, 4'd4, 16'd76};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 76, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4901] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4902] = {5'd0, 4'd8, 4'd0, 16'd67};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 67, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4903] = {5'd1, 4'd2, 4'd4, 16'd77};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 77, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4904] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4905] = {5'd0, 4'd8, 4'd0, 16'd111};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 111, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4906] = {5'd1, 4'd2, 4'd4, 16'd78};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 78, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4907] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4908] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4909] = {5'd1, 4'd2, 4'd4, 16'd79};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 79, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4910] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4911] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4912] = {5'd1, 4'd2, 4'd4, 16'd80};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 80, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4913] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4914] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4915] = {5'd1, 4'd2, 4'd4, 16'd81};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 81, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4916] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4917] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4918] = {5'd1, 4'd2, 4'd4, 16'd82};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 82, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4919] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4920] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4921] = {5'd1, 4'd2, 4'd4, 16'd83};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 83, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4922] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4923] = {5'd0, 4'd8, 4'd0, 16'd45};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 45, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4924] = {5'd1, 4'd2, 4'd4, 16'd84};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 84, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4925] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4926] = {5'd0, 4'd8, 4'd0, 16'd84};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 84, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4927] = {5'd1, 4'd2, 4'd4, 16'd85};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 85, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4928] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4929] = {5'd0, 4'd8, 4'd0, 16'd121};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 121, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4930] = {5'd1, 4'd2, 4'd4, 16'd86};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 86, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4931] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4932] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4933] = {5'd1, 4'd2, 4'd4, 16'd87};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 87, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4934] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4935] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4936] = {5'd1, 4'd2, 4'd4, 16'd88};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 88, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4937] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4938] = {5'd0, 4'd8, 4'd0, 16'd58};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 58, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4939] = {5'd1, 4'd2, 4'd4, 16'd89};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 89, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4940] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4941] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4942] = {5'd1, 4'd2, 4'd4, 16'd90};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 90, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4943] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4944] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4945] = {5'd1, 4'd2, 4'd4, 16'd91};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 91, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4946] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4947] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4948] = {5'd1, 4'd2, 4'd4, 16'd92};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 92, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4949] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4950] = {5'd0, 4'd8, 4'd0, 16'd120};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 120, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4951] = {5'd1, 4'd2, 4'd4, 16'd93};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 93, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4952] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4953] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4954] = {5'd1, 4'd2, 4'd4, 16'd94};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 94, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4955] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4956] = {5'd0, 4'd8, 4'd0, 16'd47};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 47, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4957] = {5'd1, 4'd2, 4'd4, 16'd95};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 95, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4958] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4959] = {5'd0, 4'd8, 4'd0, 16'd104};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 104, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4960] = {5'd1, 4'd2, 4'd4, 16'd96};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 96, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4961] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4962] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4963] = {5'd1, 4'd2, 4'd4, 16'd97};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 97, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4964] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4965] = {5'd0, 4'd8, 4'd0, 16'd109};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 109, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4966] = {5'd1, 4'd2, 4'd4, 16'd98};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 98, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4967] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4968] = {5'd0, 4'd8, 4'd0, 16'd108};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 108, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4969] = {5'd1, 4'd2, 4'd4, 16'd99};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 99, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4970] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4971] = {5'd0, 4'd8, 4'd0, 16'd13};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 13, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4972] = {5'd1, 4'd2, 4'd4, 16'd100};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 100, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4973] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4974] = {5'd0, 4'd8, 4'd0, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 10, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4975] = {5'd1, 4'd2, 4'd4, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 101, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4976] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4977] = {5'd0, 4'd8, 4'd0, 16'd67};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 67, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4978] = {5'd1, 4'd2, 4'd4, 16'd102};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 102, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4979] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4980] = {5'd0, 4'd8, 4'd0, 16'd111};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 111, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4981] = {5'd1, 4'd2, 4'd4, 16'd103};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 103, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4982] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4983] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4984] = {5'd1, 4'd2, 4'd4, 16'd104};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 104, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4985] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4986] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4987] = {5'd1, 4'd2, 4'd4, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 105, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4988] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4989] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4990] = {5'd1, 4'd2, 4'd4, 16'd106};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 106, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4991] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4992] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4993] = {5'd1, 4'd2, 4'd4, 16'd107};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 107, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4994] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4995] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4996] = {5'd1, 4'd2, 4'd4, 16'd108};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 108, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[4997] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[4998] = {5'd0, 4'd8, 4'd0, 16'd45};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 45, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[4999] = {5'd1, 4'd2, 4'd4, 16'd109};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 109, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[5000] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[5001] = {5'd0, 4'd8, 4'd0, 16'd76};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 76, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[5002] = {5'd1, 4'd2, 4'd4, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 110, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[5003] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[5004] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[5005] = {5'd1, 4'd2, 4'd4, 16'd111};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 111, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[5006] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[5007] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[5008] = {5'd1, 4'd2, 4'd4, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 112, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[5009] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[5010] = {5'd0, 4'd8, 4'd0, 16'd103};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 103, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[5011] = {5'd1, 4'd2, 4'd4, 16'd113};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 113, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[5012] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[5013] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[5014] = {5'd1, 4'd2, 4'd4, 16'd114};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 114, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[5015] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[5016] = {5'd0, 4'd8, 4'd0, 16'd104};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 104, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[5017] = {5'd1, 4'd2, 4'd4, 16'd115};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 115, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[5018] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[5019] = {5'd0, 4'd8, 4'd0, 16'd58};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 58, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[5020] = {5'd1, 4'd2, 4'd4, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 116, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[5021] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[5022] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[5023] = {5'd1, 4'd2, 4'd4, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 117, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[5024] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[5025] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'literal'}
    instructions[5026] = {5'd1, 4'd2, 4'd4, 16'd118};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 4, 'literal': 118, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'addl'}
    instructions[5027] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 111, 'op': 'store'}
    instructions[5028] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 118 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 118, 'op': 'literal'}
    instructions[5029] = {5'd1, 4'd2, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 118 {'a': 4, 'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 118, 'op': 'addl'}
    instructions[5030] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 118 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 118, 'op': 'store'}
    instructions[5031] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119, 'op': 'addl'}
    instructions[5032] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119, 'op': 'addl'}
    instructions[5033] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119, 'op': 'load'}
    instructions[5034] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119, 'op': 'store'}
    instructions[5035] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119, 'op': 'addl'}
    instructions[5036] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119, 'op': 'addl'}
    instructions[5037] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119, 'op': 'addl'}
    instructions[5038] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119, 'op': 'load'}
    instructions[5039] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5040] = {5'd5, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119, 'op': 'load'}
    instructions[5041] = {5'd11, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119, 'op': 'add'}
    instructions[5042] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119, 'op': 'addl'}
    instructions[5043] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119, 'op': 'load'}
    instructions[5044] = {5'd8, 4'd0, 4'd8, 16'd5064};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 121 {'a': 8, 'label': 5064, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 121, 'op': 'jmp_if_false'}
    instructions[5045] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119, 'op': 'addl'}
    instructions[5046] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119, 'op': 'addl'}
    instructions[5047] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119, 'op': 'load'}
    instructions[5048] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119, 'op': 'store'}
    instructions[5049] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119, 'op': 'addl'}
    instructions[5050] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119, 'op': 'literal'}
    instructions[5051] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119, 'op': 'store'}
    instructions[5052] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119, 'op': 'addl'}
    instructions[5053] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119, 'op': 'addl'}
    instructions[5054] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119, 'op': 'addl'}
    instructions[5055] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119, 'op': 'load'}
    instructions[5056] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5057] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119, 'op': 'load'}
    instructions[5058] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119, 'op': 'add'}
    instructions[5059] = {5'd1, 4'd2, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119 {'a': 4, 'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119, 'op': 'addl'}
    instructions[5060] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119, 'op': 'store'}
    instructions[5061] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5062] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119, 'op': 'load'}
    instructions[5063] = {5'd12, 4'd0, 4'd0, 16'd5065};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 121 {'label': 5065, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 121, 'op': 'goto'}
    instructions[5064] = {5'd12, 4'd0, 4'd0, 16'd5066};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 121 {'label': 5066, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 121, 'op': 'goto'}
    instructions[5065] = {5'd12, 4'd0, 4'd0, 16'd5031};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119 {'label': 5031, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 119, 'op': 'goto'}
    instructions[5066] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 121 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 121, 'op': 'literal'}
    instructions[5067] = {5'd1, 4'd2, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 121 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 121, 'op': 'addl'}
    instructions[5068] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 121 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 121, 'op': 'store'}
    instructions[5069] = {5'd1, 4'd8, 4'd4, 16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122 {'a': 4, 'literal': 5, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122, 'op': 'addl'}
    instructions[5070] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122, 'op': 'store'}
    instructions[5071] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122, 'op': 'addl'}
    instructions[5072] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122, 'op': 'addl'}
    instructions[5073] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122, 'op': 'addl'}
    instructions[5074] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122, 'op': 'load'}
    instructions[5075] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5076] = {5'd5, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122, 'op': 'load'}
    instructions[5077] = {5'd11, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122, 'op': 'add'}
    instructions[5078] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122, 'op': 'addl'}
    instructions[5079] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122, 'op': 'load'}
    instructions[5080] = {5'd8, 4'd0, 4'd8, 16'd5100};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 125 {'a': 8, 'label': 5100, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 125, 'op': 'jmp_if_false'}
    instructions[5081] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122, 'op': 'addl'}
    instructions[5082] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122, 'op': 'addl'}
    instructions[5083] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122, 'op': 'load'}
    instructions[5084] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122, 'op': 'store'}
    instructions[5085] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122, 'op': 'addl'}
    instructions[5086] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122, 'op': 'literal'}
    instructions[5087] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122, 'op': 'store'}
    instructions[5088] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122, 'op': 'addl'}
    instructions[5089] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122, 'op': 'addl'}
    instructions[5090] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122, 'op': 'addl'}
    instructions[5091] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122, 'op': 'load'}
    instructions[5092] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5093] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122, 'op': 'load'}
    instructions[5094] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122, 'op': 'add'}
    instructions[5095] = {5'd1, 4'd2, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122, 'op': 'addl'}
    instructions[5096] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122, 'op': 'store'}
    instructions[5097] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5098] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122, 'op': 'load'}
    instructions[5099] = {5'd12, 4'd0, 4'd0, 16'd5101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 125 {'label': 5101, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 125, 'op': 'goto'}
    instructions[5100] = {5'd12, 4'd0, 4'd0, 16'd5102};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 125 {'label': 5102, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 125, 'op': 'goto'}
    instructions[5101] = {5'd12, 4'd0, 4'd0, 16'd5069};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122 {'label': 5069, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 122, 'op': 'goto'}
    instructions[5102] = {5'd0, 4'd8, 4'd0, 16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 125 {'literal': 5, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 125, 'op': 'literal'}
    instructions[5103] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 125 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 125, 'op': 'store'}
    instructions[5104] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 125 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 125, 'op': 'addl'}
    instructions[5105] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 125 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 125, 'op': 'addl'}
    instructions[5106] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 125 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 125, 'op': 'addl'}
    instructions[5107] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 125 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 125, 'op': 'load'}
    instructions[5108] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 125 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 125, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5109] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 125 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 125, 'op': 'load'}
    instructions[5110] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 125 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 125, 'op': 'add'}
    instructions[5111] = {5'd1, 4'd2, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 125 {'a': 4, 'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 125, 'op': 'addl'}
    instructions[5112] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 125 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 125, 'op': 'store'}
    instructions[5113] = {5'd0, 4'd8, 4'd0, 16'd9};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127 {'literal': 9, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127, 'op': 'literal'}
    instructions[5114] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127, 'op': 'store'}
    instructions[5115] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127, 'op': 'addl'}
    instructions[5116] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127, 'op': 'addl'}
    instructions[5117] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127, 'op': 'addl'}
    instructions[5118] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127, 'op': 'load'}
    instructions[5119] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5120] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127, 'op': 'load'}
    instructions[5121] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127, 'op': 'unsigned_greater'}
    instructions[5122] = {5'd8, 4'd0, 4'd8, 16'd5142};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127 {'a': 8, 'label': 5142, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127, 'op': 'jmp_if_false'}
    instructions[5123] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127, 'op': 'addl'}
    instructions[5124] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127, 'op': 'addl'}
    instructions[5125] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127, 'op': 'load'}
    instructions[5126] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127, 'op': 'store'}
    instructions[5127] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127, 'op': 'addl'}
    instructions[5128] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127, 'op': 'literal'}
    instructions[5129] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127, 'op': 'store'}
    instructions[5130] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127, 'op': 'addl'}
    instructions[5131] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127, 'op': 'addl'}
    instructions[5132] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127, 'op': 'addl'}
    instructions[5133] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127, 'op': 'load'}
    instructions[5134] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5135] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127, 'op': 'load'}
    instructions[5136] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127, 'op': 'add'}
    instructions[5137] = {5'd1, 4'd2, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127 {'a': 4, 'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127, 'op': 'addl'}
    instructions[5138] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127, 'op': 'store'}
    instructions[5139] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5140] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127, 'op': 'load'}
    instructions[5141] = {5'd12, 4'd0, 4'd0, 16'd5142};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127 {'label': 5142, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 127, 'op': 'goto'}
    instructions[5142] = {5'd0, 4'd8, 4'd0, 16'd99};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128 {'literal': 99, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128, 'op': 'literal'}
    instructions[5143] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128, 'op': 'store'}
    instructions[5144] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128, 'op': 'addl'}
    instructions[5145] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128, 'op': 'addl'}
    instructions[5146] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128, 'op': 'addl'}
    instructions[5147] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128, 'op': 'load'}
    instructions[5148] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5149] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128, 'op': 'load'}
    instructions[5150] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128, 'op': 'unsigned_greater'}
    instructions[5151] = {5'd8, 4'd0, 4'd8, 16'd5171};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128 {'a': 8, 'label': 5171, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128, 'op': 'jmp_if_false'}
    instructions[5152] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128, 'op': 'addl'}
    instructions[5153] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128, 'op': 'addl'}
    instructions[5154] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128, 'op': 'load'}
    instructions[5155] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128, 'op': 'store'}
    instructions[5156] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128, 'op': 'addl'}
    instructions[5157] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128, 'op': 'literal'}
    instructions[5158] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128, 'op': 'store'}
    instructions[5159] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128, 'op': 'addl'}
    instructions[5160] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128, 'op': 'addl'}
    instructions[5161] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128, 'op': 'addl'}
    instructions[5162] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128, 'op': 'load'}
    instructions[5163] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5164] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128, 'op': 'load'}
    instructions[5165] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128, 'op': 'add'}
    instructions[5166] = {5'd1, 4'd2, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128 {'a': 4, 'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128, 'op': 'addl'}
    instructions[5167] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128, 'op': 'store'}
    instructions[5168] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5169] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128, 'op': 'load'}
    instructions[5170] = {5'd12, 4'd0, 4'd0, 16'd5171};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128 {'label': 5171, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 128, 'op': 'goto'}
    instructions[5171] = {5'd0, 4'd8, 4'd0, 16'd999};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129 {'literal': 999, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129, 'op': 'literal'}
    instructions[5172] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129, 'op': 'store'}
    instructions[5173] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129, 'op': 'addl'}
    instructions[5174] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129, 'op': 'addl'}
    instructions[5175] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129, 'op': 'addl'}
    instructions[5176] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129, 'op': 'load'}
    instructions[5177] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5178] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129, 'op': 'load'}
    instructions[5179] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129, 'op': 'unsigned_greater'}
    instructions[5180] = {5'd8, 4'd0, 4'd8, 16'd5200};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129 {'a': 8, 'label': 5200, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129, 'op': 'jmp_if_false'}
    instructions[5181] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129, 'op': 'addl'}
    instructions[5182] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129, 'op': 'addl'}
    instructions[5183] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129, 'op': 'load'}
    instructions[5184] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129, 'op': 'store'}
    instructions[5185] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129, 'op': 'addl'}
    instructions[5186] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129, 'op': 'literal'}
    instructions[5187] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129, 'op': 'store'}
    instructions[5188] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129, 'op': 'addl'}
    instructions[5189] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129, 'op': 'addl'}
    instructions[5190] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129, 'op': 'addl'}
    instructions[5191] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129, 'op': 'load'}
    instructions[5192] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5193] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129, 'op': 'load'}
    instructions[5194] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129, 'op': 'add'}
    instructions[5195] = {5'd1, 4'd2, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129 {'a': 4, 'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129, 'op': 'addl'}
    instructions[5196] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129, 'op': 'store'}
    instructions[5197] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5198] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129, 'op': 'load'}
    instructions[5199] = {5'd12, 4'd0, 4'd0, 16'd5200};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129 {'label': 5200, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 129, 'op': 'goto'}
    instructions[5200] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 131 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 131, 'op': 'store'}
    instructions[5201] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 131 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 131, 'op': 'addl'}
    instructions[5202] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 131 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 131, 'op': 'store'}
    instructions[5203] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 131 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 131, 'op': 'addl'}
    instructions[5204] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 131 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 131, 'op': 'addl'}
    instructions[5205] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 131 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 131, 'op': 'addl'}
    instructions[5206] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 131 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 131, 'op': 'load'}
    instructions[5207] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 131 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 131, 'op': 'store'}
    instructions[5208] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 131 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 131, 'op': 'addl'}
    instructions[5209] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 131 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 131, 'op': 'addl'}
    instructions[5210] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 131 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 131, 'op': 'addl'}
    instructions[5211] = {5'd3, 4'd6, 4'd0, 16'd5537};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 131 {'z': 6, 'label': 5537, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 131, 'op': 'call'}
    instructions[5212] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 131 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 131, 'op': 'addl'}
    instructions[5213] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 131 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 131, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5214] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 131 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 131, 'op': 'load'}
    instructions[5215] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 131 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 131, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5216] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 131 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 131, 'op': 'load'}
    instructions[5217] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 131 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 131, 'op': 'addl'}
    instructions[5218] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 133 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 133, 'op': 'store'}
    instructions[5219] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 133 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 133, 'op': 'addl'}
    instructions[5220] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 133 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 133, 'op': 'store'}
    instructions[5221] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 133 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 133, 'op': 'addl'}
    instructions[5222] = {5'd1, 4'd8, 4'd4, 16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 133 {'a': 4, 'literal': 5, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 133, 'op': 'addl'}
    instructions[5223] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 133 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 133, 'op': 'store'}
    instructions[5224] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 133 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 133, 'op': 'addl'}
    instructions[5225] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 133 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 133, 'op': 'addl'}
    instructions[5226] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 133 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 133, 'op': 'addl'}
    instructions[5227] = {5'd3, 4'd6, 4'd0, 16'd5553};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 133 {'z': 6, 'label': 5553, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 133, 'op': 'call'}
    instructions[5228] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 133 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 133, 'op': 'addl'}
    instructions[5229] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 133 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 133, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5230] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 133 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 133, 'op': 'load'}
    instructions[5231] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 133 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 133, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5232] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 133 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 133, 'op': 'load'}
    instructions[5233] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 133 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 133, 'op': 'addl'}
    instructions[5234] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 134 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 134, 'op': 'store'}
    instructions[5235] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 134 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 134, 'op': 'addl'}
    instructions[5236] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 134 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 134, 'op': 'store'}
    instructions[5237] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 134 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 134, 'op': 'addl'}
    instructions[5238] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 134 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 134, 'op': 'addl'}
    instructions[5239] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 134 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 134, 'op': 'addl'}
    instructions[5240] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 134 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 134, 'op': 'load'}
    instructions[5241] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 134 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 134, 'op': 'store'}
    instructions[5242] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 134 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 134, 'op': 'addl'}
    instructions[5243] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 134 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 134, 'op': 'addl'}
    instructions[5244] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 134 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 134, 'op': 'addl'}
    instructions[5245] = {5'd3, 4'd6, 4'd0, 16'd5720};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 134 {'z': 6, 'label': 5720, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 134, 'op': 'call'}
    instructions[5246] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 134 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 134, 'op': 'addl'}
    instructions[5247] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 134 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 134, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5248] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 134 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 134, 'op': 'load'}
    instructions[5249] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 134 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 134, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5250] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 134 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 134, 'op': 'load'}
    instructions[5251] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 134 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 134, 'op': 'addl'}
    instructions[5252] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135, 'op': 'store'}
    instructions[5253] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135, 'op': 'addl'}
    instructions[5254] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135, 'op': 'store'}
    instructions[5255] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135, 'op': 'addl'}
    instructions[5256] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135, 'op': 'literal'}
    instructions[5257] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135, 'op': 'store'}
    instructions[5258] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135, 'op': 'addl'}
    instructions[5259] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135, 'op': 'addl'}
    instructions[5260] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135, 'op': 'addl'}
    instructions[5261] = {5'd3, 4'd6, 4'd0, 16'd5553};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135 {'z': 6, 'label': 5553, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135, 'op': 'call'}
    instructions[5262] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135, 'op': 'addl'}
    instructions[5263] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5264] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135, 'op': 'load'}
    instructions[5265] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5266] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135, 'op': 'load'}
    instructions[5267] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 135, 'op': 'addl'}
    instructions[5268] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 136 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 136, 'op': 'store'}
    instructions[5269] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 136 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 136, 'op': 'addl'}
    instructions[5270] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 136 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 136, 'op': 'store'}
    instructions[5271] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 136 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 136, 'op': 'addl'}
    instructions[5272] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 136 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 136, 'op': 'addl'}
    instructions[5273] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 136 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 136, 'op': 'addl'}
    instructions[5274] = {5'd3, 4'd6, 4'd0, 16'd6136};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 136 {'z': 6, 'label': 6136, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 136, 'op': 'call'}
    instructions[5275] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 136 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 136, 'op': 'addl'}
    instructions[5276] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 136 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 136, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5277] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 136 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 136, 'op': 'load'}
    instructions[5278] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 136 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 136, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5279] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 136 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 136, 'op': 'load'}
    instructions[5280] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 136 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 136, 'op': 'addl'}
    instructions[5281] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 138 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 138, 'op': 'addl'}
    instructions[5282] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 138 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 138, 'op': 'addl'}
    instructions[5283] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 138 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 138, 'op': 'load'}
    instructions[5284] = {5'd1, 4'd2, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 138 {'a': 4, 'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 138, 'op': 'addl'}
    instructions[5285] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 138 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 138, 'op': 'store'}
    instructions[5286] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 139 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 139, 'op': 'literal'}
    instructions[5287] = {5'd1, 4'd2, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 139 {'a': 4, 'literal': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 139, 'op': 'addl'}
    instructions[5288] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 139 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 139, 'op': 'store'}
    instructions[5289] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 140 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 140, 'op': 'literal'}
    instructions[5290] = {5'd1, 4'd2, 4'd4, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 140 {'a': 4, 'literal': 4, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 140, 'op': 'addl'}
    instructions[5291] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 140 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 140, 'op': 'store'}
    instructions[5292] = {5'd0, 4'd8, 4'd0, 16'd1046};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 141 {'literal': 1046, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 141, 'op': 'literal'}
    instructions[5293] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 141 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 141, 'op': 'store'}
    instructions[5294] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 141 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 141, 'op': 'addl'}
    instructions[5295] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 141 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 141, 'op': 'addl'}
    instructions[5296] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 141 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 141, 'op': 'addl'}
    instructions[5297] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 141 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 141, 'op': 'load'}
    instructions[5298] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 141 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 141, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5299] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 141 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 141, 'op': 'load'}
    instructions[5300] = {5'd20, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 141 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 141, 'op': 'unsigned_greater_equal'}
    instructions[5301] = {5'd8, 4'd0, 4'd8, 16'd5421};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 150 {'a': 8, 'label': 5421, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 150, 'op': 'jmp_if_false'}
    instructions[5302] = {5'd0, 4'd8, 4'd0, 16'd1046};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 142 {'literal': 1046, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 142, 'op': 'literal'}
    instructions[5303] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 142 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 142, 'op': 'store'}
    instructions[5304] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 142 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 142, 'op': 'addl'}
    instructions[5305] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 142 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 142, 'op': 'addl'}
    instructions[5306] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 142 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 142, 'op': 'addl'}
    instructions[5307] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 142 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 142, 'op': 'load'}
    instructions[5308] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 142 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 142, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5309] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 142 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 142, 'op': 'load'}
    instructions[5310] = {5'd21, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 142 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 142, 'op': 'subtract'}
    instructions[5311] = {5'd1, 4'd2, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 142 {'a': 4, 'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 142, 'op': 'addl'}
    instructions[5312] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 142 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 142, 'op': 'store'}
    instructions[5313] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 143 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 143, 'op': 'store'}
    instructions[5314] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 143 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 143, 'op': 'addl'}
    instructions[5315] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 143 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 143, 'op': 'store'}
    instructions[5316] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 143 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 143, 'op': 'addl'}
    instructions[5317] = {5'd0, 4'd8, 4'd0, 16'd1046};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 143 {'literal': 1046, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 143, 'op': 'literal'}
    instructions[5318] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 143 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 143, 'op': 'store'}
    instructions[5319] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 143 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 143, 'op': 'addl'}
    instructions[5320] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 143 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 143, 'op': 'addl'}
    instructions[5321] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 143 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 143, 'op': 'addl'}
    instructions[5322] = {5'd3, 4'd6, 4'd0, 16'd5537};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 143 {'z': 6, 'label': 5537, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 143, 'op': 'call'}
    instructions[5323] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 143 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 143, 'op': 'addl'}
    instructions[5324] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 143 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 143, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5325] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 143 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 143, 'op': 'load'}
    instructions[5326] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 143 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 143, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5327] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 143 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 143, 'op': 'load'}
    instructions[5328] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 143 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 143, 'op': 'addl'}
    instructions[5329] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144, 'op': 'literal'}
    instructions[5330] = {5'd1, 4'd2, 4'd4, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144 {'a': 4, 'literal': 4, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144, 'op': 'addl'}
    instructions[5331] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144, 'op': 'store'}
    instructions[5332] = {5'd1, 4'd8, 4'd4, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144 {'a': 4, 'literal': 4, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144, 'op': 'addl'}
    instructions[5333] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144, 'op': 'addl'}
    instructions[5334] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144, 'op': 'load'}
    instructions[5335] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144, 'op': 'store'}
    instructions[5336] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144, 'op': 'addl'}
    instructions[5337] = {5'd0, 4'd8, 4'd0, 16'd1046};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144 {'literal': 1046, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144, 'op': 'literal'}
    instructions[5338] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5339] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144, 'op': 'load'}
    instructions[5340] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144, 'op': 'unsigned_greater'}
    instructions[5341] = {5'd8, 4'd0, 4'd8, 16'd5407};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144 {'a': 8, 'label': 5407, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144, 'op': 'jmp_if_false'}
    instructions[5342] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145, 'op': 'store'}
    instructions[5343] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145, 'op': 'addl'}
    instructions[5344] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145, 'op': 'store'}
    instructions[5345] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145, 'op': 'addl'}
    instructions[5346] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145, 'op': 'addl'}
    instructions[5347] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145, 'op': 'addl'}
    instructions[5348] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145, 'op': 'load'}
    instructions[5349] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145, 'op': 'store'}
    instructions[5350] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145, 'op': 'addl'}
    instructions[5351] = {5'd1, 4'd8, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145 {'a': 4, 'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145, 'op': 'addl'}
    instructions[5352] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145, 'op': 'addl'}
    instructions[5353] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145, 'op': 'load'}
    instructions[5354] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5355] = {5'd5, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145, 'op': 'load'}
    instructions[5356] = {5'd11, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145, 'op': 'add'}
    instructions[5357] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145, 'op': 'addl'}
    instructions[5358] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145, 'op': 'load'}
    instructions[5359] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145, 'op': 'store'}
    instructions[5360] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145, 'op': 'addl'}
    instructions[5361] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145, 'op': 'addl'}
    instructions[5362] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145, 'op': 'addl'}
    instructions[5363] = {5'd3, 4'd6, 4'd0, 16'd5623};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145 {'z': 6, 'label': 5623, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145, 'op': 'call'}
    instructions[5364] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145, 'op': 'addl'}
    instructions[5365] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5366] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145, 'op': 'load'}
    instructions[5367] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5368] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145, 'op': 'load'}
    instructions[5369] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 145, 'op': 'addl'}
    instructions[5370] = {5'd1, 4'd8, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 146 {'a': 4, 'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 146, 'op': 'addl'}
    instructions[5371] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 146 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 146, 'op': 'addl'}
    instructions[5372] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 146 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 146, 'op': 'load'}
    instructions[5373] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 146 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 146, 'op': 'store'}
    instructions[5374] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 146 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 146, 'op': 'addl'}
    instructions[5375] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 146 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 146, 'op': 'literal'}
    instructions[5376] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 146 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 146, 'op': 'store'}
    instructions[5377] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 146 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 146, 'op': 'addl'}
    instructions[5378] = {5'd1, 4'd8, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 146 {'a': 4, 'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 146, 'op': 'addl'}
    instructions[5379] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 146 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 146, 'op': 'addl'}
    instructions[5380] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 146 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 146, 'op': 'load'}
    instructions[5381] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 146 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 146, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5382] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 146 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 146, 'op': 'load'}
    instructions[5383] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 146 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 146, 'op': 'add'}
    instructions[5384] = {5'd1, 4'd2, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 146 {'a': 4, 'literal': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 146, 'op': 'addl'}
    instructions[5385] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 146 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 146, 'op': 'store'}
    instructions[5386] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 146 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 146, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5387] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 146 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 146, 'op': 'load'}
    instructions[5388] = {5'd1, 4'd8, 4'd4, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144 {'a': 4, 'literal': 4, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144, 'op': 'addl'}
    instructions[5389] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144, 'op': 'addl'}
    instructions[5390] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144, 'op': 'load'}
    instructions[5391] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144, 'op': 'store'}
    instructions[5392] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144, 'op': 'addl'}
    instructions[5393] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144, 'op': 'literal'}
    instructions[5394] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144, 'op': 'store'}
    instructions[5395] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144, 'op': 'addl'}
    instructions[5396] = {5'd1, 4'd8, 4'd4, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144 {'a': 4, 'literal': 4, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144, 'op': 'addl'}
    instructions[5397] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144, 'op': 'addl'}
    instructions[5398] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144, 'op': 'load'}
    instructions[5399] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5400] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144, 'op': 'load'}
    instructions[5401] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144, 'op': 'add'}
    instructions[5402] = {5'd1, 4'd2, 4'd4, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144 {'a': 4, 'literal': 4, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144, 'op': 'addl'}
    instructions[5403] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144, 'op': 'store'}
    instructions[5404] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5405] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144, 'op': 'load'}
    instructions[5406] = {5'd12, 4'd0, 4'd0, 16'd5332};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144 {'label': 5332, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 144, 'op': 'goto'}
    instructions[5407] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 148 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 148, 'op': 'store'}
    instructions[5408] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 148 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 148, 'op': 'addl'}
    instructions[5409] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 148 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 148, 'op': 'store'}
    instructions[5410] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 148 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 148, 'op': 'addl'}
    instructions[5411] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 148 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 148, 'op': 'addl'}
    instructions[5412] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 148 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 148, 'op': 'addl'}
    instructions[5413] = {5'd3, 4'd6, 4'd0, 16'd6136};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 148 {'z': 6, 'label': 6136, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 148, 'op': 'call'}
    instructions[5414] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 148 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 148, 'op': 'addl'}
    instructions[5415] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 148 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 148, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5416] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 148 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 148, 'op': 'load'}
    instructions[5417] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 148 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 148, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5418] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 148 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 148, 'op': 'load'}
    instructions[5419] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 148 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 148, 'op': 'addl'}
    instructions[5420] = {5'd12, 4'd0, 4'd0, 16'd5422};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 150 {'label': 5422, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 150, 'op': 'goto'}
    instructions[5421] = {5'd12, 4'd0, 4'd0, 16'd5423};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 150 {'label': 5423, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 150, 'op': 'goto'}
    instructions[5422] = {5'd12, 4'd0, 4'd0, 16'd5292};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 141 {'label': 5292, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 141, 'op': 'goto'}
    instructions[5423] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 150 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 150, 'op': 'store'}
    instructions[5424] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 150 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 150, 'op': 'addl'}
    instructions[5425] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 150 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 150, 'op': 'store'}
    instructions[5426] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 150 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 150, 'op': 'addl'}
    instructions[5427] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 150 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 150, 'op': 'addl'}
    instructions[5428] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 150 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 150, 'op': 'addl'}
    instructions[5429] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 150 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 150, 'op': 'load'}
    instructions[5430] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 150 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 150, 'op': 'store'}
    instructions[5431] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 150 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 150, 'op': 'addl'}
    instructions[5432] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 150 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 150, 'op': 'addl'}
    instructions[5433] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 150 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 150, 'op': 'addl'}
    instructions[5434] = {5'd3, 4'd6, 4'd0, 16'd5537};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 150 {'z': 6, 'label': 5537, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 150, 'op': 'call'}
    instructions[5435] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 150 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 150, 'op': 'addl'}
    instructions[5436] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 150 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 150, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5437] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 150 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 150, 'op': 'load'}
    instructions[5438] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 150 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 150, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5439] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 150 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 150, 'op': 'load'}
    instructions[5440] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 150 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 150, 'op': 'addl'}
    instructions[5441] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151, 'op': 'literal'}
    instructions[5442] = {5'd1, 4'd2, 4'd4, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151 {'a': 4, 'literal': 4, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151, 'op': 'addl'}
    instructions[5443] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151, 'op': 'store'}
    instructions[5444] = {5'd1, 4'd8, 4'd4, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151 {'a': 4, 'literal': 4, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151, 'op': 'addl'}
    instructions[5445] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151, 'op': 'addl'}
    instructions[5446] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151, 'op': 'load'}
    instructions[5447] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151, 'op': 'store'}
    instructions[5448] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151, 'op': 'addl'}
    instructions[5449] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151, 'op': 'addl'}
    instructions[5450] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151, 'op': 'addl'}
    instructions[5451] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151, 'op': 'load'}
    instructions[5452] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5453] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151, 'op': 'load'}
    instructions[5454] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151, 'op': 'unsigned_greater'}
    instructions[5455] = {5'd8, 4'd0, 4'd8, 16'd5521};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151 {'a': 8, 'label': 5521, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151, 'op': 'jmp_if_false'}
    instructions[5456] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152, 'op': 'store'}
    instructions[5457] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152, 'op': 'addl'}
    instructions[5458] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152, 'op': 'store'}
    instructions[5459] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152, 'op': 'addl'}
    instructions[5460] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152, 'op': 'addl'}
    instructions[5461] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152, 'op': 'addl'}
    instructions[5462] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152, 'op': 'load'}
    instructions[5463] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152, 'op': 'store'}
    instructions[5464] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152, 'op': 'addl'}
    instructions[5465] = {5'd1, 4'd8, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152 {'a': 4, 'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152, 'op': 'addl'}
    instructions[5466] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152, 'op': 'addl'}
    instructions[5467] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152, 'op': 'load'}
    instructions[5468] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5469] = {5'd5, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152, 'op': 'load'}
    instructions[5470] = {5'd11, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152, 'op': 'add'}
    instructions[5471] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152, 'op': 'addl'}
    instructions[5472] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152, 'op': 'load'}
    instructions[5473] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152, 'op': 'store'}
    instructions[5474] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152, 'op': 'addl'}
    instructions[5475] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152, 'op': 'addl'}
    instructions[5476] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152, 'op': 'addl'}
    instructions[5477] = {5'd3, 4'd6, 4'd0, 16'd5623};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152 {'z': 6, 'label': 5623, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152, 'op': 'call'}
    instructions[5478] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152, 'op': 'addl'}
    instructions[5479] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5480] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152, 'op': 'load'}
    instructions[5481] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5482] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152, 'op': 'load'}
    instructions[5483] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 152, 'op': 'addl'}
    instructions[5484] = {5'd1, 4'd8, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 153 {'a': 4, 'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 153, 'op': 'addl'}
    instructions[5485] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 153 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 153, 'op': 'addl'}
    instructions[5486] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 153 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 153, 'op': 'load'}
    instructions[5487] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 153 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 153, 'op': 'store'}
    instructions[5488] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 153 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 153, 'op': 'addl'}
    instructions[5489] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 153 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 153, 'op': 'literal'}
    instructions[5490] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 153 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 153, 'op': 'store'}
    instructions[5491] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 153 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 153, 'op': 'addl'}
    instructions[5492] = {5'd1, 4'd8, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 153 {'a': 4, 'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 153, 'op': 'addl'}
    instructions[5493] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 153 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 153, 'op': 'addl'}
    instructions[5494] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 153 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 153, 'op': 'load'}
    instructions[5495] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 153 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 153, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5496] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 153 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 153, 'op': 'load'}
    instructions[5497] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 153 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 153, 'op': 'add'}
    instructions[5498] = {5'd1, 4'd2, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 153 {'a': 4, 'literal': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 153, 'op': 'addl'}
    instructions[5499] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 153 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 153, 'op': 'store'}
    instructions[5500] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 153 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 153, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5501] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 153 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 153, 'op': 'load'}
    instructions[5502] = {5'd1, 4'd8, 4'd4, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151 {'a': 4, 'literal': 4, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151, 'op': 'addl'}
    instructions[5503] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151, 'op': 'addl'}
    instructions[5504] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151, 'op': 'load'}
    instructions[5505] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151, 'op': 'store'}
    instructions[5506] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151, 'op': 'addl'}
    instructions[5507] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151, 'op': 'literal'}
    instructions[5508] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151, 'op': 'store'}
    instructions[5509] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151, 'op': 'addl'}
    instructions[5510] = {5'd1, 4'd8, 4'd4, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151 {'a': 4, 'literal': 4, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151, 'op': 'addl'}
    instructions[5511] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151, 'op': 'addl'}
    instructions[5512] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151, 'op': 'load'}
    instructions[5513] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5514] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151, 'op': 'load'}
    instructions[5515] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151, 'op': 'add'}
    instructions[5516] = {5'd1, 4'd2, 4'd4, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151 {'a': 4, 'literal': 4, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151, 'op': 'addl'}
    instructions[5517] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151, 'op': 'store'}
    instructions[5518] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5519] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151, 'op': 'load'}
    instructions[5520] = {5'd12, 4'd0, 4'd0, 16'd5444};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151 {'label': 5444, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 151, 'op': 'goto'}
    instructions[5521] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 155 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 155, 'op': 'store'}
    instructions[5522] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 155 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 155, 'op': 'addl'}
    instructions[5523] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 155 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 155, 'op': 'store'}
    instructions[5524] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 155 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 155, 'op': 'addl'}
    instructions[5525] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 155 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 155, 'op': 'addl'}
    instructions[5526] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 155 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 155, 'op': 'addl'}
    instructions[5527] = {5'd3, 4'd6, 4'd0, 16'd6136};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 155 {'z': 6, 'label': 6136, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 155, 'op': 'call'}
    instructions[5528] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 155 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 155, 'op': 'addl'}
    instructions[5529] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 155 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 155, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5530] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 155 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 155, 'op': 'load'}
    instructions[5531] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 155 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 155, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5532] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 155 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 155, 'op': 'load'}
    instructions[5533] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 155 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 155, 'op': 'addl'}
    instructions[5534] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 106 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 106, 'op': 'addl'}
    instructions[5535] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 106 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 106, 'op': 'addl'}
    instructions[5536] = {5'd19, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 106 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 106, 'op': 'return'}
    instructions[5537] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 30 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 30, 'op': 'addl'}
    instructions[5538] = {5'd0, 4'd8, 4'd0, 16'd95};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 31 {'literal': 95, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 31, 'op': 'literal'}
    instructions[5539] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 31 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 31, 'op': 'addl'}
    instructions[5540] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 31 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 31, 'op': 'load'}
    instructions[5541] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 31 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 31, 'op': 'store'}
    instructions[5542] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 31 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 31, 'op': 'addl'}
    instructions[5543] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 31 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 31, 'op': 'addl'}
    instructions[5544] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 31 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 31, 'op': 'addl'}
    instructions[5545] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 31 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 31, 'op': 'load'}
    instructions[5546] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 31 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 31, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5547] = {5'd5, 4'd0, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 31 {'a': 3, 'z': 0, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 31, 'op': 'load'}
    instructions[5548] = {5'd17, 4'd0, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 31 {'a': 0, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 31, 'op': 'write'}
    instructions[5549] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 31 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 31, 'op': 'addl'}
    instructions[5550] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 30 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 30, 'op': 'addl'}
    instructions[5551] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 30 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 30, 'op': 'addl'}
    instructions[5552] = {5'd19, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 30 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/application.c : 30, 'op': 'return'}
    instructions[5553] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 34 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 34, 'op': 'addl'}
    instructions[5554] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 35 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 35, 'op': 'literal'}
    instructions[5555] = {5'd1, 4'd2, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 35 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 35, 'op': 'addl'}
    instructions[5556] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 35 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 35, 'op': 'store'}
    instructions[5557] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 36 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 36, 'op': 'addl'}
    instructions[5558] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 36 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 36, 'op': 'addl'}
    instructions[5559] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 36 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 36, 'op': 'load'}
    instructions[5560] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 36 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 36, 'op': 'store'}
    instructions[5561] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 36 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 36, 'op': 'addl'}
    instructions[5562] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 36 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 36, 'op': 'addl'}
    instructions[5563] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 36 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 36, 'op': 'addl'}
    instructions[5564] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 36 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 36, 'op': 'load'}
    instructions[5565] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 36 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 36, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5566] = {5'd5, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 36 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 36, 'op': 'load'}
    instructions[5567] = {5'd11, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 36 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 36, 'op': 'add'}
    instructions[5568] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 36 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 36, 'op': 'addl'}
    instructions[5569] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 36 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 36, 'op': 'load'}
    instructions[5570] = {5'd8, 4'd0, 4'd8, 16'd5618};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 40 {'a': 8, 'label': 5618, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 40, 'op': 'jmp_if_false'}
    instructions[5571] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37, 'op': 'store'}
    instructions[5572] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37, 'op': 'addl'}
    instructions[5573] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37, 'op': 'store'}
    instructions[5574] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37, 'op': 'addl'}
    instructions[5575] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37, 'op': 'addl'}
    instructions[5576] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37, 'op': 'addl'}
    instructions[5577] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37, 'op': 'load'}
    instructions[5578] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37, 'op': 'store'}
    instructions[5579] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37, 'op': 'addl'}
    instructions[5580] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37, 'op': 'addl'}
    instructions[5581] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37, 'op': 'addl'}
    instructions[5582] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37, 'op': 'load'}
    instructions[5583] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5584] = {5'd5, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37, 'op': 'load'}
    instructions[5585] = {5'd11, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37, 'op': 'add'}
    instructions[5586] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37, 'op': 'addl'}
    instructions[5587] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37, 'op': 'load'}
    instructions[5588] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37, 'op': 'store'}
    instructions[5589] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37, 'op': 'addl'}
    instructions[5590] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37, 'op': 'addl'}
    instructions[5591] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37, 'op': 'addl'}
    instructions[5592] = {5'd3, 4'd6, 4'd0, 16'd5623};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37 {'z': 6, 'label': 5623, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37, 'op': 'call'}
    instructions[5593] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37, 'op': 'addl'}
    instructions[5594] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5595] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37, 'op': 'load'}
    instructions[5596] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5597] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37, 'op': 'load'}
    instructions[5598] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 37, 'op': 'addl'}
    instructions[5599] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 38 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 38, 'op': 'addl'}
    instructions[5600] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 38 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 38, 'op': 'addl'}
    instructions[5601] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 38 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 38, 'op': 'load'}
    instructions[5602] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 38 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 38, 'op': 'store'}
    instructions[5603] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 38 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 38, 'op': 'addl'}
    instructions[5604] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 38 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 38, 'op': 'literal'}
    instructions[5605] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 38 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 38, 'op': 'store'}
    instructions[5606] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 38 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 38, 'op': 'addl'}
    instructions[5607] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 38 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 38, 'op': 'addl'}
    instructions[5608] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 38 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 38, 'op': 'addl'}
    instructions[5609] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 38 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 38, 'op': 'load'}
    instructions[5610] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 38 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 38, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5611] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 38 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 38, 'op': 'load'}
    instructions[5612] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 38 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 38, 'op': 'add'}
    instructions[5613] = {5'd1, 4'd2, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 38 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 38, 'op': 'addl'}
    instructions[5614] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 38 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 38, 'op': 'store'}
    instructions[5615] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 38 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 38, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5616] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 38 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 38, 'op': 'load'}
    instructions[5617] = {5'd12, 4'd0, 4'd0, 16'd5619};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 40 {'label': 5619, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 40, 'op': 'goto'}
    instructions[5618] = {5'd12, 4'd0, 4'd0, 16'd5620};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 40 {'label': 5620, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 40, 'op': 'goto'}
    instructions[5619] = {5'd12, 4'd0, 4'd0, 16'd5557};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 36 {'label': 5557, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 36, 'op': 'goto'}
    instructions[5620] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 34 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 34, 'op': 'addl'}
    instructions[5621] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 34 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 34, 'op': 'addl'}
    instructions[5622] = {5'd19, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 34 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 34, 'op': 'return'}
    instructions[5623] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 17 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 17, 'op': 'addl'}
    instructions[5624] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 18 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 18, 'op': 'store'}
    instructions[5625] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 18 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 18, 'op': 'addl'}
    instructions[5626] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 18 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 18, 'op': 'store'}
    instructions[5627] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 18 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 18, 'op': 'addl'}
    instructions[5628] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 18 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 18, 'op': 'addl'}
    instructions[5629] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 18 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 18, 'op': 'addl'}
    instructions[5630] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 18 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 18, 'op': 'load'}
    instructions[5631] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 18 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 18, 'op': 'store'}
    instructions[5632] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 18 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 18, 'op': 'addl'}
    instructions[5633] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 18 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 18, 'op': 'addl'}
    instructions[5634] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 18 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 18, 'op': 'addl'}
    instructions[5635] = {5'd3, 4'd6, 4'd0, 16'd5704};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 18 {'z': 6, 'label': 5704, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 18, 'op': 'call'}
    instructions[5636] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 18 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 18, 'op': 'addl'}
    instructions[5637] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 18 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 18, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5638] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 18 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 18, 'op': 'load'}
    instructions[5639] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 18 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 18, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5640] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 18 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 18, 'op': 'load'}
    instructions[5641] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 18 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 18, 'op': 'addl'}
    instructions[5642] = {5'd0, 4'd8, 4'd0, 16'd51};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 19 {'literal': 51, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 19, 'op': 'literal'}
    instructions[5643] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 19 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 19, 'op': 'addl'}
    instructions[5644] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 19 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 19, 'op': 'load'}
    instructions[5645] = {5'd8, 4'd0, 4'd8, 16'd5661};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 19 {'a': 8, 'label': 5661, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 19, 'op': 'jmp_if_false'}
    instructions[5646] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 20 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 20, 'op': 'literal'}
    instructions[5647] = {5'd0, 4'd2, 4'd0, 16'd51};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 20 {'literal': 51, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 20, 'op': 'literal'}
    instructions[5648] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 20 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 20, 'op': 'store'}
    instructions[5649] = {5'd0, 4'd8, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 21 {'literal': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 21, 'op': 'literal'}
    instructions[5650] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 21 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 21, 'op': 'store'}
    instructions[5651] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 21 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 21, 'op': 'addl'}
    instructions[5652] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 21 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 21, 'op': 'addl'}
    instructions[5653] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 21 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 21, 'op': 'addl'}
    instructions[5654] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 21 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 21, 'op': 'load'}
    instructions[5655] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 21 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 21, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5656] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 21 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 21, 'op': 'load'}
    instructions[5657] = {5'd22, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 21 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 21, 'op': 'shift_left'}
    instructions[5658] = {5'd0, 4'd2, 4'd0, 16'd53};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 21 {'literal': 53, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 21, 'op': 'literal'}
    instructions[5659] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 21 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 21, 'op': 'store'}
    instructions[5660] = {5'd12, 4'd0, 4'd0, 16'd5701};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 19 {'label': 5701, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 19, 'op': 'goto'}
    instructions[5661] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 23 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 23, 'op': 'literal'}
    instructions[5662] = {5'd0, 4'd2, 4'd0, 16'd51};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 23 {'literal': 51, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 23, 'op': 'literal'}
    instructions[5663] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 23 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 23, 'op': 'store'}
    instructions[5664] = {5'd0, 4'd8, 4'd0, 16'd255};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 24 {'literal': 255, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 24, 'op': 'literal'}
    instructions[5665] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 24 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 24, 'op': 'store'}
    instructions[5666] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 24 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 24, 'op': 'addl'}
    instructions[5667] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 24 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 24, 'op': 'addl'}
    instructions[5668] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 24 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 24, 'op': 'addl'}
    instructions[5669] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 24 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 24, 'op': 'load'}
    instructions[5670] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 24 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 24, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5671] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 24 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 24, 'op': 'load'}
    instructions[5672] = {5'd10, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 24 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 24, 'op': 'and'}
    instructions[5673] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 24 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 24, 'op': 'store'}
    instructions[5674] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 24 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 24, 'op': 'addl'}
    instructions[5675] = {5'd0, 4'd8, 4'd0, 16'd53};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 24 {'literal': 53, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 24, 'op': 'literal'}
    instructions[5676] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 24 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 24, 'op': 'addl'}
    instructions[5677] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 24 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 24, 'op': 'load'}
    instructions[5678] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 24 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 24, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5679] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 24 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 24, 'op': 'load'}
    instructions[5680] = {5'd16, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 24 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 24, 'op': 'or'}
    instructions[5681] = {5'd0, 4'd2, 4'd0, 16'd53};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 24 {'literal': 53, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 24, 'op': 'literal'}
    instructions[5682] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 24 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 24, 'op': 'store'}
    instructions[5683] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 25 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 25, 'op': 'store'}
    instructions[5684] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 25 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 25, 'op': 'addl'}
    instructions[5685] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 25 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 25, 'op': 'store'}
    instructions[5686] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 25 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 25, 'op': 'addl'}
    instructions[5687] = {5'd0, 4'd8, 4'd0, 16'd53};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 25 {'literal': 53, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 25, 'op': 'literal'}
    instructions[5688] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 25 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 25, 'op': 'addl'}
    instructions[5689] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 25 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 25, 'op': 'load'}
    instructions[5690] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 25 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 25, 'op': 'store'}
    instructions[5691] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 25 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 25, 'op': 'addl'}
    instructions[5692] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 25 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 25, 'op': 'addl'}
    instructions[5693] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 25 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 25, 'op': 'addl'}
    instructions[5694] = {5'd3, 4'd6, 4'd0, 16'd5537};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 25 {'z': 6, 'label': 5537, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 25, 'op': 'call'}
    instructions[5695] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 25 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 25, 'op': 'addl'}
    instructions[5696] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 25 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 25, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5697] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 25 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 25, 'op': 'load'}
    instructions[5698] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 25 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 25, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5699] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 25 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 25, 'op': 'load'}
    instructions[5700] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 25 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 25, 'op': 'addl'}
    instructions[5701] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 17 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 17, 'op': 'addl'}
    instructions[5702] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 17 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 17, 'op': 'addl'}
    instructions[5703] = {5'd19, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 17 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 17, 'op': 'return'}
    instructions[5704] = {5'd1, 4'd3, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 95 {'a': 3, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 95, 'op': 'addl'}
    instructions[5705] = {5'd0, 4'd8, 4'd0, 16'd7};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 96 {'literal': 7, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 96, 'op': 'literal'}
    instructions[5706] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 96 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 96, 'op': 'addl'}
    instructions[5707] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 96 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 96, 'op': 'load'}
    instructions[5708] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 96 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 96, 'op': 'store'}
    instructions[5709] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 96 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 96, 'op': 'addl'}
    instructions[5710] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 96 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 96, 'op': 'addl'}
    instructions[5711] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 96 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 96, 'op': 'addl'}
    instructions[5712] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 96 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 96, 'op': 'load'}
    instructions[5713] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 96 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 96, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5714] = {5'd5, 4'd0, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 96 {'a': 3, 'z': 0, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 96, 'op': 'load'}
    instructions[5715] = {5'd17, 4'd0, 4'd0, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 96 {'a': 0, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 96, 'op': 'write'}
    instructions[5716] = {5'd1, 4'd3, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 96 {'a': 3, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 96, 'op': 'addl'}
    instructions[5717] = {5'd1, 4'd3, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 95 {'a': 4, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 95, 'op': 'addl'}
    instructions[5718] = {5'd1, 4'd4, 4'd7, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 95 {'a': 7, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 95, 'op': 'addl'}
    instructions[5719] = {5'd19, 4'd0, 4'd6, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 95 {'a': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 95, 'op': 'return'}
    instructions[5720] = {5'd1, 4'd3, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 42 {'a': 3, 'literal': 6, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 42, 'op': 'addl'}
    instructions[5721] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 43 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 43, 'op': 'literal'}
    instructions[5722] = {5'd1, 4'd2, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 43 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 43, 'op': 'addl'}
    instructions[5723] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 43 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 43, 'op': 'store'}
    instructions[5724] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 44 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 44, 'op': 'literal'}
    instructions[5725] = {5'd1, 4'd2, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 44 {'a': 4, 'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 44, 'op': 'addl'}
    instructions[5726] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 44 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 44, 'op': 'store'}
    instructions[5727] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 45 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 45, 'op': 'literal'}
    instructions[5728] = {5'd1, 4'd2, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 45 {'a': 4, 'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 45, 'op': 'addl'}
    instructions[5729] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 45 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 45, 'op': 'store'}
    instructions[5730] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 46 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 46, 'op': 'literal'}
    instructions[5731] = {5'd1, 4'd2, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 46 {'a': 4, 'literal': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 46, 'op': 'addl'}
    instructions[5732] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 46 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 46, 'op': 'store'}
    instructions[5733] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 47 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 47, 'op': 'literal'}
    instructions[5734] = {5'd1, 4'd2, 4'd4, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 47 {'a': 4, 'literal': 4, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 47, 'op': 'addl'}
    instructions[5735] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 47 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 47, 'op': 'store'}
    instructions[5736] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 48 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 48, 'op': 'literal'}
    instructions[5737] = {5'd1, 4'd2, 4'd4, 16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 48 {'a': 4, 'literal': 5, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 48, 'op': 'addl'}
    instructions[5738] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 48 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 48, 'op': 'store'}
    instructions[5739] = {5'd0, 4'd8, 4'd0, 16'd10000};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 50 {'literal': 10000, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 50, 'op': 'literal'}
    instructions[5740] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 50 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 50, 'op': 'store'}
    instructions[5741] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 50 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 50, 'op': 'addl'}
    instructions[5742] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 50 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 50, 'op': 'addl'}
    instructions[5743] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 50 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 50, 'op': 'addl'}
    instructions[5744] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 50 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 50, 'op': 'load'}
    instructions[5745] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 50 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 50, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5746] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 50 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 50, 'op': 'load'}
    instructions[5747] = {5'd20, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 50 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 50, 'op': 'unsigned_greater_equal'}
    instructions[5748] = {5'd8, 4'd0, 4'd8, 16'd5779};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 54 {'a': 8, 'label': 5779, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 54, 'op': 'jmp_if_false'}
    instructions[5749] = {5'd1, 4'd8, 4'd4, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 51 {'a': 4, 'literal': 4, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 51, 'op': 'addl'}
    instructions[5750] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 51 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 51, 'op': 'addl'}
    instructions[5751] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 51 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 51, 'op': 'load'}
    instructions[5752] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 51 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 51, 'op': 'store'}
    instructions[5753] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 51 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 51, 'op': 'addl'}
    instructions[5754] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 51 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 51, 'op': 'literal'}
    instructions[5755] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 51 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 51, 'op': 'store'}
    instructions[5756] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 51 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 51, 'op': 'addl'}
    instructions[5757] = {5'd1, 4'd8, 4'd4, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 51 {'a': 4, 'literal': 4, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 51, 'op': 'addl'}
    instructions[5758] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 51 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 51, 'op': 'addl'}
    instructions[5759] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 51 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 51, 'op': 'load'}
    instructions[5760] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 51 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 51, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5761] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 51 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 51, 'op': 'load'}
    instructions[5762] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 51 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 51, 'op': 'add'}
    instructions[5763] = {5'd1, 4'd2, 4'd4, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 51 {'a': 4, 'literal': 4, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 51, 'op': 'addl'}
    instructions[5764] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 51 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 51, 'op': 'store'}
    instructions[5765] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 51 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 51, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5766] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 51 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 51, 'op': 'load'}
    instructions[5767] = {5'd0, 4'd8, 4'd0, 16'd10000};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 52 {'literal': 10000, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 52, 'op': 'literal'}
    instructions[5768] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 52 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 52, 'op': 'store'}
    instructions[5769] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 52 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 52, 'op': 'addl'}
    instructions[5770] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 52 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 52, 'op': 'addl'}
    instructions[5771] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 52 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 52, 'op': 'addl'}
    instructions[5772] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 52 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 52, 'op': 'load'}
    instructions[5773] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 52 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 52, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5774] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 52 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 52, 'op': 'load'}
    instructions[5775] = {5'd21, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 52 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 52, 'op': 'subtract'}
    instructions[5776] = {5'd1, 4'd2, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 52 {'a': 4, 'literal': -1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 52, 'op': 'addl'}
    instructions[5777] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 52 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 52, 'op': 'store'}
    instructions[5778] = {5'd12, 4'd0, 4'd0, 16'd5780};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 54 {'label': 5780, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 54, 'op': 'goto'}
    instructions[5779] = {5'd12, 4'd0, 4'd0, 16'd5781};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 54 {'label': 5781, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 54, 'op': 'goto'}
    instructions[5780] = {5'd12, 4'd0, 4'd0, 16'd5739};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 50 {'label': 5739, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 50, 'op': 'goto'}
    instructions[5781] = {5'd1, 4'd8, 4'd4, 16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 54 {'a': 4, 'literal': 5, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 54, 'op': 'addl'}
    instructions[5782] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 54 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 54, 'op': 'addl'}
    instructions[5783] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 54 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 54, 'op': 'load'}
    instructions[5784] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 54 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 54, 'op': 'store'}
    instructions[5785] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 54 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 54, 'op': 'addl'}
    instructions[5786] = {5'd1, 4'd8, 4'd4, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 54 {'a': 4, 'literal': 4, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 54, 'op': 'addl'}
    instructions[5787] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 54 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 54, 'op': 'addl'}
    instructions[5788] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 54 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 54, 'op': 'load'}
    instructions[5789] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 54 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 54, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5790] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 54 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 54, 'op': 'load'}
    instructions[5791] = {5'd16, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 54 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 54, 'op': 'or'}
    instructions[5792] = {5'd8, 4'd0, 4'd8, 16'd5821};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 54 {'a': 8, 'label': 5821, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 54, 'op': 'jmp_if_false'}
    instructions[5793] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55, 'op': 'store'}
    instructions[5794] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55, 'op': 'addl'}
    instructions[5795] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55, 'op': 'store'}
    instructions[5796] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55, 'op': 'addl'}
    instructions[5797] = {5'd1, 4'd8, 4'd4, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55 {'a': 4, 'literal': 4, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55, 'op': 'addl'}
    instructions[5798] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55, 'op': 'addl'}
    instructions[5799] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55, 'op': 'load'}
    instructions[5800] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55, 'op': 'store'}
    instructions[5801] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55, 'op': 'addl'}
    instructions[5802] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55, 'op': 'literal'}
    instructions[5803] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5804] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55, 'op': 'load'}
    instructions[5805] = {5'd16, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55, 'op': 'or'}
    instructions[5806] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55, 'op': 'store'}
    instructions[5807] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55, 'op': 'addl'}
    instructions[5808] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55, 'op': 'addl'}
    instructions[5809] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55, 'op': 'addl'}
    instructions[5810] = {5'd3, 4'd6, 4'd0, 16'd5623};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55 {'z': 6, 'label': 5623, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55, 'op': 'call'}
    instructions[5811] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55, 'op': 'addl'}
    instructions[5812] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5813] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55, 'op': 'load'}
    instructions[5814] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5815] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55, 'op': 'load'}
    instructions[5816] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 55, 'op': 'addl'}
    instructions[5817] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 56 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 56, 'op': 'literal'}
    instructions[5818] = {5'd1, 4'd2, 4'd4, 16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 56 {'a': 4, 'literal': 5, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 56, 'op': 'addl'}
    instructions[5819] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 56 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 56, 'op': 'store'}
    instructions[5820] = {5'd12, 4'd0, 4'd0, 16'd5821};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 54 {'label': 5821, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 54, 'op': 'goto'}
    instructions[5821] = {5'd0, 4'd8, 4'd0, 16'd1000};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 58 {'literal': 1000, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 58, 'op': 'literal'}
    instructions[5822] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 58 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 58, 'op': 'store'}
    instructions[5823] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 58 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 58, 'op': 'addl'}
    instructions[5824] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 58 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 58, 'op': 'addl'}
    instructions[5825] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 58 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 58, 'op': 'addl'}
    instructions[5826] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 58 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 58, 'op': 'load'}
    instructions[5827] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 58 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 58, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5828] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 58 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 58, 'op': 'load'}
    instructions[5829] = {5'd20, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 58 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 58, 'op': 'unsigned_greater_equal'}
    instructions[5830] = {5'd8, 4'd0, 4'd8, 16'd5861};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 62 {'a': 8, 'label': 5861, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 62, 'op': 'jmp_if_false'}
    instructions[5831] = {5'd1, 4'd8, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 59 {'a': 4, 'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 59, 'op': 'addl'}
    instructions[5832] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 59 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 59, 'op': 'addl'}
    instructions[5833] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 59 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 59, 'op': 'load'}
    instructions[5834] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 59 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 59, 'op': 'store'}
    instructions[5835] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 59 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 59, 'op': 'addl'}
    instructions[5836] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 59 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 59, 'op': 'literal'}
    instructions[5837] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 59 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 59, 'op': 'store'}
    instructions[5838] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 59 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 59, 'op': 'addl'}
    instructions[5839] = {5'd1, 4'd8, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 59 {'a': 4, 'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 59, 'op': 'addl'}
    instructions[5840] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 59 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 59, 'op': 'addl'}
    instructions[5841] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 59 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 59, 'op': 'load'}
    instructions[5842] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 59 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 59, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5843] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 59 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 59, 'op': 'load'}
    instructions[5844] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 59 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 59, 'op': 'add'}
    instructions[5845] = {5'd1, 4'd2, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 59 {'a': 4, 'literal': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 59, 'op': 'addl'}
    instructions[5846] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 59 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 59, 'op': 'store'}
    instructions[5847] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 59 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 59, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5848] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 59 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 59, 'op': 'load'}
    instructions[5849] = {5'd0, 4'd8, 4'd0, 16'd1000};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 60 {'literal': 1000, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 60, 'op': 'literal'}
    instructions[5850] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 60 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 60, 'op': 'store'}
    instructions[5851] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 60 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 60, 'op': 'addl'}
    instructions[5852] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 60 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 60, 'op': 'addl'}
    instructions[5853] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 60 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 60, 'op': 'addl'}
    instructions[5854] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 60 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 60, 'op': 'load'}
    instructions[5855] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 60 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 60, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5856] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 60 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 60, 'op': 'load'}
    instructions[5857] = {5'd21, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 60 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 60, 'op': 'subtract'}
    instructions[5858] = {5'd1, 4'd2, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 60 {'a': 4, 'literal': -1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 60, 'op': 'addl'}
    instructions[5859] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 60 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 60, 'op': 'store'}
    instructions[5860] = {5'd12, 4'd0, 4'd0, 16'd5862};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 62 {'label': 5862, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 62, 'op': 'goto'}
    instructions[5861] = {5'd12, 4'd0, 4'd0, 16'd5863};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 62 {'label': 5863, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 62, 'op': 'goto'}
    instructions[5862] = {5'd12, 4'd0, 4'd0, 16'd5821};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 58 {'label': 5821, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 58, 'op': 'goto'}
    instructions[5863] = {5'd1, 4'd8, 4'd4, 16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 62 {'a': 4, 'literal': 5, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 62, 'op': 'addl'}
    instructions[5864] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 62 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 62, 'op': 'addl'}
    instructions[5865] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 62 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 62, 'op': 'load'}
    instructions[5866] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 62 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 62, 'op': 'store'}
    instructions[5867] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 62 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 62, 'op': 'addl'}
    instructions[5868] = {5'd1, 4'd8, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 62 {'a': 4, 'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 62, 'op': 'addl'}
    instructions[5869] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 62 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 62, 'op': 'addl'}
    instructions[5870] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 62 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 62, 'op': 'load'}
    instructions[5871] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 62 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 62, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5872] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 62 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 62, 'op': 'load'}
    instructions[5873] = {5'd16, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 62 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 62, 'op': 'or'}
    instructions[5874] = {5'd8, 4'd0, 4'd8, 16'd5903};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 62 {'a': 8, 'label': 5903, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 62, 'op': 'jmp_if_false'}
    instructions[5875] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63, 'op': 'store'}
    instructions[5876] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63, 'op': 'addl'}
    instructions[5877] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63, 'op': 'store'}
    instructions[5878] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63, 'op': 'addl'}
    instructions[5879] = {5'd1, 4'd8, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63 {'a': 4, 'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63, 'op': 'addl'}
    instructions[5880] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63, 'op': 'addl'}
    instructions[5881] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63, 'op': 'load'}
    instructions[5882] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63, 'op': 'store'}
    instructions[5883] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63, 'op': 'addl'}
    instructions[5884] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63, 'op': 'literal'}
    instructions[5885] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5886] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63, 'op': 'load'}
    instructions[5887] = {5'd16, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63, 'op': 'or'}
    instructions[5888] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63, 'op': 'store'}
    instructions[5889] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63, 'op': 'addl'}
    instructions[5890] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63, 'op': 'addl'}
    instructions[5891] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63, 'op': 'addl'}
    instructions[5892] = {5'd3, 4'd6, 4'd0, 16'd5623};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63 {'z': 6, 'label': 5623, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63, 'op': 'call'}
    instructions[5893] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63, 'op': 'addl'}
    instructions[5894] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5895] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63, 'op': 'load'}
    instructions[5896] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5897] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63, 'op': 'load'}
    instructions[5898] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 63, 'op': 'addl'}
    instructions[5899] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 64 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 64, 'op': 'literal'}
    instructions[5900] = {5'd1, 4'd2, 4'd4, 16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 64 {'a': 4, 'literal': 5, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 64, 'op': 'addl'}
    instructions[5901] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 64 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 64, 'op': 'store'}
    instructions[5902] = {5'd12, 4'd0, 4'd0, 16'd5903};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 62 {'label': 5903, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 62, 'op': 'goto'}
    instructions[5903] = {5'd0, 4'd8, 4'd0, 16'd100};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 66 {'literal': 100, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 66, 'op': 'literal'}
    instructions[5904] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 66 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 66, 'op': 'store'}
    instructions[5905] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 66 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 66, 'op': 'addl'}
    instructions[5906] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 66 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 66, 'op': 'addl'}
    instructions[5907] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 66 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 66, 'op': 'addl'}
    instructions[5908] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 66 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 66, 'op': 'load'}
    instructions[5909] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 66 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 66, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5910] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 66 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 66, 'op': 'load'}
    instructions[5911] = {5'd20, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 66 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 66, 'op': 'unsigned_greater_equal'}
    instructions[5912] = {5'd8, 4'd0, 4'd8, 16'd5943};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 70 {'a': 8, 'label': 5943, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 70, 'op': 'jmp_if_false'}
    instructions[5913] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 67 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 67, 'op': 'addl'}
    instructions[5914] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 67 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 67, 'op': 'addl'}
    instructions[5915] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 67 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 67, 'op': 'load'}
    instructions[5916] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 67 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 67, 'op': 'store'}
    instructions[5917] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 67 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 67, 'op': 'addl'}
    instructions[5918] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 67 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 67, 'op': 'literal'}
    instructions[5919] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 67 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 67, 'op': 'store'}
    instructions[5920] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 67 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 67, 'op': 'addl'}
    instructions[5921] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 67 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 67, 'op': 'addl'}
    instructions[5922] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 67 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 67, 'op': 'addl'}
    instructions[5923] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 67 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 67, 'op': 'load'}
    instructions[5924] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 67 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 67, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5925] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 67 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 67, 'op': 'load'}
    instructions[5926] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 67 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 67, 'op': 'add'}
    instructions[5927] = {5'd1, 4'd2, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 67 {'a': 4, 'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 67, 'op': 'addl'}
    instructions[5928] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 67 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 67, 'op': 'store'}
    instructions[5929] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 67 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 67, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5930] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 67 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 67, 'op': 'load'}
    instructions[5931] = {5'd0, 4'd8, 4'd0, 16'd100};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 68 {'literal': 100, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 68, 'op': 'literal'}
    instructions[5932] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 68 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 68, 'op': 'store'}
    instructions[5933] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 68 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 68, 'op': 'addl'}
    instructions[5934] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 68 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 68, 'op': 'addl'}
    instructions[5935] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 68 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 68, 'op': 'addl'}
    instructions[5936] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 68 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 68, 'op': 'load'}
    instructions[5937] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 68 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 68, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5938] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 68 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 68, 'op': 'load'}
    instructions[5939] = {5'd21, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 68 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 68, 'op': 'subtract'}
    instructions[5940] = {5'd1, 4'd2, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 68 {'a': 4, 'literal': -1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 68, 'op': 'addl'}
    instructions[5941] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 68 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 68, 'op': 'store'}
    instructions[5942] = {5'd12, 4'd0, 4'd0, 16'd5944};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 70 {'label': 5944, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 70, 'op': 'goto'}
    instructions[5943] = {5'd12, 4'd0, 4'd0, 16'd5945};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 70 {'label': 5945, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 70, 'op': 'goto'}
    instructions[5944] = {5'd12, 4'd0, 4'd0, 16'd5903};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 66 {'label': 5903, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 66, 'op': 'goto'}
    instructions[5945] = {5'd1, 4'd8, 4'd4, 16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 70 {'a': 4, 'literal': 5, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 70, 'op': 'addl'}
    instructions[5946] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 70 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 70, 'op': 'addl'}
    instructions[5947] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 70 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 70, 'op': 'load'}
    instructions[5948] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 70 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 70, 'op': 'store'}
    instructions[5949] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 70 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 70, 'op': 'addl'}
    instructions[5950] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 70 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 70, 'op': 'addl'}
    instructions[5951] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 70 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 70, 'op': 'addl'}
    instructions[5952] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 70 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 70, 'op': 'load'}
    instructions[5953] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 70 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 70, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5954] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 70 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 70, 'op': 'load'}
    instructions[5955] = {5'd16, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 70 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 70, 'op': 'or'}
    instructions[5956] = {5'd8, 4'd0, 4'd8, 16'd5985};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 70 {'a': 8, 'label': 5985, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 70, 'op': 'jmp_if_false'}
    instructions[5957] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71, 'op': 'store'}
    instructions[5958] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71, 'op': 'addl'}
    instructions[5959] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71, 'op': 'store'}
    instructions[5960] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71, 'op': 'addl'}
    instructions[5961] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71, 'op': 'addl'}
    instructions[5962] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71, 'op': 'addl'}
    instructions[5963] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71, 'op': 'load'}
    instructions[5964] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71, 'op': 'store'}
    instructions[5965] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71, 'op': 'addl'}
    instructions[5966] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71, 'op': 'literal'}
    instructions[5967] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5968] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71, 'op': 'load'}
    instructions[5969] = {5'd16, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71, 'op': 'or'}
    instructions[5970] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71, 'op': 'store'}
    instructions[5971] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71, 'op': 'addl'}
    instructions[5972] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71, 'op': 'addl'}
    instructions[5973] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71, 'op': 'addl'}
    instructions[5974] = {5'd3, 4'd6, 4'd0, 16'd5623};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71 {'z': 6, 'label': 5623, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71, 'op': 'call'}
    instructions[5975] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71, 'op': 'addl'}
    instructions[5976] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5977] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71, 'op': 'load'}
    instructions[5978] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5979] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71, 'op': 'load'}
    instructions[5980] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 71, 'op': 'addl'}
    instructions[5981] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 72 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 72, 'op': 'literal'}
    instructions[5982] = {5'd1, 4'd2, 4'd4, 16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 72 {'a': 4, 'literal': 5, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 72, 'op': 'addl'}
    instructions[5983] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 72 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 72, 'op': 'store'}
    instructions[5984] = {5'd12, 4'd0, 4'd0, 16'd5985};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 70 {'label': 5985, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 70, 'op': 'goto'}
    instructions[5985] = {5'd0, 4'd8, 4'd0, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 74 {'literal': 10, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 74, 'op': 'literal'}
    instructions[5986] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 74 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 74, 'op': 'store'}
    instructions[5987] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 74 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 74, 'op': 'addl'}
    instructions[5988] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 74 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 74, 'op': 'addl'}
    instructions[5989] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 74 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 74, 'op': 'addl'}
    instructions[5990] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 74 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 74, 'op': 'load'}
    instructions[5991] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 74 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 74, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5992] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 74 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 74, 'op': 'load'}
    instructions[5993] = {5'd20, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 74 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 74, 'op': 'unsigned_greater_equal'}
    instructions[5994] = {5'd8, 4'd0, 4'd8, 16'd6025};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 78 {'a': 8, 'label': 6025, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 78, 'op': 'jmp_if_false'}
    instructions[5995] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 75 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 75, 'op': 'addl'}
    instructions[5996] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 75 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 75, 'op': 'addl'}
    instructions[5997] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 75 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 75, 'op': 'load'}
    instructions[5998] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 75 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 75, 'op': 'store'}
    instructions[5999] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 75 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 75, 'op': 'addl'}
    instructions[6000] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 75 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 75, 'op': 'literal'}
    instructions[6001] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 75 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 75, 'op': 'store'}
    instructions[6002] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 75 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 75, 'op': 'addl'}
    instructions[6003] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 75 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 75, 'op': 'addl'}
    instructions[6004] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 75 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 75, 'op': 'addl'}
    instructions[6005] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 75 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 75, 'op': 'load'}
    instructions[6006] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 75 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 75, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[6007] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 75 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 75, 'op': 'load'}
    instructions[6008] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 75 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 75, 'op': 'add'}
    instructions[6009] = {5'd1, 4'd2, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 75 {'a': 4, 'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 75, 'op': 'addl'}
    instructions[6010] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 75 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 75, 'op': 'store'}
    instructions[6011] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 75 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 75, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[6012] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 75 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 75, 'op': 'load'}
    instructions[6013] = {5'd0, 4'd8, 4'd0, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 76 {'literal': 10, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 76, 'op': 'literal'}
    instructions[6014] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 76 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 76, 'op': 'store'}
    instructions[6015] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 76 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 76, 'op': 'addl'}
    instructions[6016] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 76 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 76, 'op': 'addl'}
    instructions[6017] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 76 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 76, 'op': 'addl'}
    instructions[6018] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 76 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 76, 'op': 'load'}
    instructions[6019] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 76 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 76, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[6020] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 76 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 76, 'op': 'load'}
    instructions[6021] = {5'd21, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 76 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 76, 'op': 'subtract'}
    instructions[6022] = {5'd1, 4'd2, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 76 {'a': 4, 'literal': -1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 76, 'op': 'addl'}
    instructions[6023] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 76 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 76, 'op': 'store'}
    instructions[6024] = {5'd12, 4'd0, 4'd0, 16'd6026};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 78 {'label': 6026, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 78, 'op': 'goto'}
    instructions[6025] = {5'd12, 4'd0, 4'd0, 16'd6027};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 78 {'label': 6027, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 78, 'op': 'goto'}
    instructions[6026] = {5'd12, 4'd0, 4'd0, 16'd5985};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 74 {'label': 5985, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 74, 'op': 'goto'}
    instructions[6027] = {5'd1, 4'd8, 4'd4, 16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 78 {'a': 4, 'literal': 5, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 78, 'op': 'addl'}
    instructions[6028] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 78 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 78, 'op': 'addl'}
    instructions[6029] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 78 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 78, 'op': 'load'}
    instructions[6030] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 78 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 78, 'op': 'store'}
    instructions[6031] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 78 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 78, 'op': 'addl'}
    instructions[6032] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 78 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 78, 'op': 'addl'}
    instructions[6033] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 78 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 78, 'op': 'addl'}
    instructions[6034] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 78 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 78, 'op': 'load'}
    instructions[6035] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 78 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 78, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[6036] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 78 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 78, 'op': 'load'}
    instructions[6037] = {5'd16, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 78 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 78, 'op': 'or'}
    instructions[6038] = {5'd8, 4'd0, 4'd8, 16'd6067};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 78 {'a': 8, 'label': 6067, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 78, 'op': 'jmp_if_false'}
    instructions[6039] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79, 'op': 'store'}
    instructions[6040] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79, 'op': 'addl'}
    instructions[6041] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79, 'op': 'store'}
    instructions[6042] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79, 'op': 'addl'}
    instructions[6043] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79, 'op': 'addl'}
    instructions[6044] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79, 'op': 'addl'}
    instructions[6045] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79, 'op': 'load'}
    instructions[6046] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79, 'op': 'store'}
    instructions[6047] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79, 'op': 'addl'}
    instructions[6048] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79, 'op': 'literal'}
    instructions[6049] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[6050] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79, 'op': 'load'}
    instructions[6051] = {5'd16, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79, 'op': 'or'}
    instructions[6052] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79, 'op': 'store'}
    instructions[6053] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79, 'op': 'addl'}
    instructions[6054] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79, 'op': 'addl'}
    instructions[6055] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79, 'op': 'addl'}
    instructions[6056] = {5'd3, 4'd6, 4'd0, 16'd5623};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79 {'z': 6, 'label': 5623, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79, 'op': 'call'}
    instructions[6057] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79, 'op': 'addl'}
    instructions[6058] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[6059] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79, 'op': 'load'}
    instructions[6060] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[6061] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79, 'op': 'load'}
    instructions[6062] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 79, 'op': 'addl'}
    instructions[6063] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 80 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 80, 'op': 'literal'}
    instructions[6064] = {5'd1, 4'd2, 4'd4, 16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 80 {'a': 4, 'literal': 5, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 80, 'op': 'addl'}
    instructions[6065] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 80 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 80, 'op': 'store'}
    instructions[6066] = {5'd12, 4'd0, 4'd0, 16'd6067};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 78 {'label': 6067, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 78, 'op': 'goto'}
    instructions[6067] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 82 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 82, 'op': 'literal'}
    instructions[6068] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 82 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 82, 'op': 'store'}
    instructions[6069] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 82 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 82, 'op': 'addl'}
    instructions[6070] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 82 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 82, 'op': 'addl'}
    instructions[6071] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 82 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 82, 'op': 'addl'}
    instructions[6072] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 82 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 82, 'op': 'load'}
    instructions[6073] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 82 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 82, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[6074] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 82 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 82, 'op': 'load'}
    instructions[6075] = {5'd20, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 82 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 82, 'op': 'unsigned_greater_equal'}
    instructions[6076] = {5'd8, 4'd0, 4'd8, 16'd6107};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86 {'a': 8, 'label': 6107, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86, 'op': 'jmp_if_false'}
    instructions[6077] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 83 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 83, 'op': 'addl'}
    instructions[6078] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 83 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 83, 'op': 'addl'}
    instructions[6079] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 83 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 83, 'op': 'load'}
    instructions[6080] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 83 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 83, 'op': 'store'}
    instructions[6081] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 83 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 83, 'op': 'addl'}
    instructions[6082] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 83 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 83, 'op': 'literal'}
    instructions[6083] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 83 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 83, 'op': 'store'}
    instructions[6084] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 83 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 83, 'op': 'addl'}
    instructions[6085] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 83 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 83, 'op': 'addl'}
    instructions[6086] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 83 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 83, 'op': 'addl'}
    instructions[6087] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 83 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 83, 'op': 'load'}
    instructions[6088] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 83 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 83, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[6089] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 83 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 83, 'op': 'load'}
    instructions[6090] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 83 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 83, 'op': 'add'}
    instructions[6091] = {5'd1, 4'd2, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 83 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 83, 'op': 'addl'}
    instructions[6092] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 83 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 83, 'op': 'store'}
    instructions[6093] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 83 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 83, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[6094] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 83 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 83, 'op': 'load'}
    instructions[6095] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 84 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 84, 'op': 'literal'}
    instructions[6096] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 84 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 84, 'op': 'store'}
    instructions[6097] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 84 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 84, 'op': 'addl'}
    instructions[6098] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 84 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 84, 'op': 'addl'}
    instructions[6099] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 84 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 84, 'op': 'addl'}
    instructions[6100] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 84 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 84, 'op': 'load'}
    instructions[6101] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 84 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 84, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[6102] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 84 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 84, 'op': 'load'}
    instructions[6103] = {5'd21, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 84 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 84, 'op': 'subtract'}
    instructions[6104] = {5'd1, 4'd2, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 84 {'a': 4, 'literal': -1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 84, 'op': 'addl'}
    instructions[6105] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 84 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 84, 'op': 'store'}
    instructions[6106] = {5'd12, 4'd0, 4'd0, 16'd6108};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86 {'label': 6108, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86, 'op': 'goto'}
    instructions[6107] = {5'd12, 4'd0, 4'd0, 16'd6109};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86 {'label': 6109, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86, 'op': 'goto'}
    instructions[6108] = {5'd12, 4'd0, 4'd0, 16'd6067};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 82 {'label': 6067, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 82, 'op': 'goto'}
    instructions[6109] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86, 'op': 'store'}
    instructions[6110] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86, 'op': 'addl'}
    instructions[6111] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86, 'op': 'store'}
    instructions[6112] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86, 'op': 'addl'}
    instructions[6113] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86, 'op': 'addl'}
    instructions[6114] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86, 'op': 'addl'}
    instructions[6115] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86, 'op': 'load'}
    instructions[6116] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86, 'op': 'store'}
    instructions[6117] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86, 'op': 'addl'}
    instructions[6118] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86, 'op': 'literal'}
    instructions[6119] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[6120] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86, 'op': 'load'}
    instructions[6121] = {5'd16, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86, 'op': 'or'}
    instructions[6122] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86, 'op': 'store'}
    instructions[6123] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86, 'op': 'addl'}
    instructions[6124] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86, 'op': 'addl'}
    instructions[6125] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86, 'op': 'addl'}
    instructions[6126] = {5'd3, 4'd6, 4'd0, 16'd5623};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86 {'z': 6, 'label': 5623, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86, 'op': 'call'}
    instructions[6127] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86, 'op': 'addl'}
    instructions[6128] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[6129] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86, 'op': 'load'}
    instructions[6130] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[6131] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86, 'op': 'load'}
    instructions[6132] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 86, 'op': 'addl'}
    instructions[6133] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 42 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 42, 'op': 'addl'}
    instructions[6134] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 42 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 42, 'op': 'addl'}
    instructions[6135] = {5'd19, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 42 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 42, 'op': 'return'}
    instructions[6136] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 29 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 29, 'op': 'addl'}
    instructions[6137] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30, 'op': 'literal'}
    instructions[6138] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30, 'op': 'store'}
    instructions[6139] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30, 'op': 'addl'}
    instructions[6140] = {5'd0, 4'd8, 4'd0, 16'd51};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30 {'literal': 51, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30, 'op': 'literal'}
    instructions[6141] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30, 'op': 'addl'}
    instructions[6142] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30, 'op': 'load'}
    instructions[6143] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[6144] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30, 'op': 'load'}
    instructions[6145] = {5'd13, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30, 'op': 'equal'}
    instructions[6146] = {5'd8, 4'd0, 4'd8, 16'd6166};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30 {'a': 8, 'label': 6166, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30, 'op': 'jmp_if_false'}
    instructions[6147] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30, 'op': 'store'}
    instructions[6148] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30, 'op': 'addl'}
    instructions[6149] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30, 'op': 'store'}
    instructions[6150] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30, 'op': 'addl'}
    instructions[6151] = {5'd0, 4'd8, 4'd0, 16'd53};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30 {'literal': 53, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30, 'op': 'literal'}
    instructions[6152] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30, 'op': 'addl'}
    instructions[6153] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30, 'op': 'load'}
    instructions[6154] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30, 'op': 'store'}
    instructions[6155] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30, 'op': 'addl'}
    instructions[6156] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30, 'op': 'addl'}
    instructions[6157] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30, 'op': 'addl'}
    instructions[6158] = {5'd3, 4'd6, 4'd0, 16'd5537};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30 {'z': 6, 'label': 5537, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30, 'op': 'call'}
    instructions[6159] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30, 'op': 'addl'}
    instructions[6160] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[6161] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30, 'op': 'load'}
    instructions[6162] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[6163] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30, 'op': 'load'}
    instructions[6164] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30, 'op': 'addl'}
    instructions[6165] = {5'd12, 4'd0, 4'd0, 16'd6166};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30 {'label': 6166, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 30, 'op': 'goto'}
    instructions[6166] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 31 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 31, 'op': 'literal'}
    instructions[6167] = {5'd0, 4'd2, 4'd0, 16'd51};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 31 {'literal': 51, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 31, 'op': 'literal'}
    instructions[6168] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 31 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 31, 'op': 'store'}
    instructions[6169] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 29 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 29, 'op': 'addl'}
    instructions[6170] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 29 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 29, 'op': 'addl'}
    instructions[6171] = {5'd19, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 29 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 29, 'op': 'return'}
    instructions[6172] = {5'd1, 4'd3, 4'd3, 16'd127};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 89 {'a': 3, 'literal': 127, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 89, 'op': 'addl'}
    instructions[6173] = {5'd0, 4'd8, 4'd0, 16'd72};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 72, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6174] = {5'd1, 4'd2, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6175] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6176] = {5'd0, 4'd8, 4'd0, 16'd84};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 84, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6177] = {5'd1, 4'd2, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6178] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6179] = {5'd0, 4'd8, 4'd0, 16'd84};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 84, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6180] = {5'd1, 4'd2, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6181] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6182] = {5'd0, 4'd8, 4'd0, 16'd80};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 80, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6183] = {5'd1, 4'd2, 4'd4, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 4, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6184] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6185] = {5'd0, 4'd8, 4'd0, 16'd47};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 47, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6186] = {5'd1, 4'd2, 4'd4, 16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 5, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6187] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6188] = {5'd0, 4'd8, 4'd0, 16'd49};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 49, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6189] = {5'd1, 4'd2, 4'd4, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 6, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6190] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6191] = {5'd0, 4'd8, 4'd0, 16'd46};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 46, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6192] = {5'd1, 4'd2, 4'd4, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 7, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6193] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6194] = {5'd0, 4'd8, 4'd0, 16'd49};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 49, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6195] = {5'd1, 4'd2, 4'd4, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 8, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6196] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6197] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6198] = {5'd1, 4'd2, 4'd4, 16'd9};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 9, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6199] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6200] = {5'd0, 4'd8, 4'd0, 16'd52};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 52, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6201] = {5'd1, 4'd2, 4'd4, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 10, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6202] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6203] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6204] = {5'd1, 4'd2, 4'd4, 16'd11};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 11, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6205] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6206] = {5'd0, 4'd8, 4'd0, 16'd52};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 52, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6207] = {5'd1, 4'd2, 4'd4, 16'd12};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 12, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6208] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6209] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6210] = {5'd1, 4'd2, 4'd4, 16'd13};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 13, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6211] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6212] = {5'd0, 4'd8, 4'd0, 16'd78};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 78, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6213] = {5'd1, 4'd2, 4'd4, 16'd14};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 14, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6214] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6215] = {5'd0, 4'd8, 4'd0, 16'd111};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 111, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6216] = {5'd1, 4'd2, 4'd4, 16'd15};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 15, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6217] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6218] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6219] = {5'd1, 4'd2, 4'd4, 16'd16};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 16, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6220] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6221] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6222] = {5'd1, 4'd2, 4'd4, 16'd17};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 17, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6223] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6224] = {5'd0, 4'd8, 4'd0, 16'd70};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 70, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6225] = {5'd1, 4'd2, 4'd4, 16'd18};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 18, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6226] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6227] = {5'd0, 4'd8, 4'd0, 16'd111};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 111, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6228] = {5'd1, 4'd2, 4'd4, 16'd19};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 19, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6229] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6230] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6231] = {5'd1, 4'd2, 4'd4, 16'd20};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 20, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6232] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6233] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6234] = {5'd1, 4'd2, 4'd4, 16'd21};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 21, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6235] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6236] = {5'd0, 4'd8, 4'd0, 16'd100};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 100, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6237] = {5'd1, 4'd2, 4'd4, 16'd22};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 22, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6238] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6239] = {5'd0, 4'd8, 4'd0, 16'd13};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 13, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6240] = {5'd1, 4'd2, 4'd4, 16'd23};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 23, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6241] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6242] = {5'd0, 4'd8, 4'd0, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 10, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6243] = {5'd1, 4'd2, 4'd4, 16'd24};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 24, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6244] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6245] = {5'd0, 4'd8, 4'd0, 16'd68};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 68, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6246] = {5'd1, 4'd2, 4'd4, 16'd25};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 25, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6247] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6248] = {5'd0, 4'd8, 4'd0, 16'd97};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 97, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6249] = {5'd1, 4'd2, 4'd4, 16'd26};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 26, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6250] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6251] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6252] = {5'd1, 4'd2, 4'd4, 16'd27};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 27, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6253] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6254] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6255] = {5'd1, 4'd2, 4'd4, 16'd28};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 28, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6256] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6257] = {5'd0, 4'd8, 4'd0, 16'd58};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 58, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6258] = {5'd1, 4'd2, 4'd4, 16'd29};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 29, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6259] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6260] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6261] = {5'd1, 4'd2, 4'd4, 16'd30};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 30, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6262] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6263] = {5'd0, 4'd8, 4'd0, 16'd84};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 84, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6264] = {5'd1, 4'd2, 4'd4, 16'd31};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 31, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6265] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6266] = {5'd0, 4'd8, 4'd0, 16'd104};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 104, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6267] = {5'd1, 4'd2, 4'd4, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 32, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6268] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6269] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6270] = {5'd1, 4'd2, 4'd4, 16'd33};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 33, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6271] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6272] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6273] = {5'd1, 4'd2, 4'd4, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 34, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6274] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6275] = {5'd0, 4'd8, 4'd0, 16'd79};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 79, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6276] = {5'd1, 4'd2, 4'd4, 16'd35};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 35, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6277] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6278] = {5'd0, 4'd8, 4'd0, 16'd99};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 99, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6279] = {5'd1, 4'd2, 4'd4, 16'd36};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 36, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6280] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6281] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6282] = {5'd1, 4'd2, 4'd4, 16'd37};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 37, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6283] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6284] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6285] = {5'd1, 4'd2, 4'd4, 16'd38};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 38, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6286] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6287] = {5'd0, 4'd8, 4'd0, 16'd51};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 51, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6288] = {5'd1, 4'd2, 4'd4, 16'd39};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 39, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6289] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6290] = {5'd0, 4'd8, 4'd0, 16'd49};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 49, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6291] = {5'd1, 4'd2, 4'd4, 16'd40};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 40, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6292] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6293] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6294] = {5'd1, 4'd2, 4'd4, 16'd41};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 41, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6295] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6296] = {5'd0, 4'd8, 4'd0, 16'd49};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 49, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6297] = {5'd1, 4'd2, 4'd4, 16'd42};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 42, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6298] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6299] = {5'd0, 4'd8, 4'd0, 16'd57};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 57, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6300] = {5'd1, 4'd2, 4'd4, 16'd43};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 43, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6301] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6302] = {5'd0, 4'd8, 4'd0, 16'd58};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 58, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6303] = {5'd1, 4'd2, 4'd4, 16'd44};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 44, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6304] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6305] = {5'd0, 4'd8, 4'd0, 16'd49};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 49, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6306] = {5'd1, 4'd2, 4'd4, 16'd45};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 45, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6307] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6308] = {5'd0, 4'd8, 4'd0, 16'd54};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 54, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6309] = {5'd1, 4'd2, 4'd4, 16'd46};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 46, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6310] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6311] = {5'd0, 4'd8, 4'd0, 16'd58};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 58, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6312] = {5'd1, 4'd2, 4'd4, 16'd47};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 47, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6313] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6314] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6315] = {5'd1, 4'd2, 4'd4, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 48, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6316] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6317] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6318] = {5'd1, 4'd2, 4'd4, 16'd49};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 49, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6319] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6320] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6321] = {5'd1, 4'd2, 4'd4, 16'd50};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 50, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6322] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6323] = {5'd0, 4'd8, 4'd0, 16'd50};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 50, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6324] = {5'd1, 4'd2, 4'd4, 16'd51};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 51, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6325] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6326] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6327] = {5'd1, 4'd2, 4'd4, 16'd52};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 52, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6328] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6329] = {5'd0, 4'd8, 4'd0, 16'd49};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 49, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6330] = {5'd1, 4'd2, 4'd4, 16'd53};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 53, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6331] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6332] = {5'd0, 4'd8, 4'd0, 16'd51};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 51, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6333] = {5'd1, 4'd2, 4'd4, 16'd54};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 54, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6334] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6335] = {5'd0, 4'd8, 4'd0, 16'd13};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 13, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6336] = {5'd1, 4'd2, 4'd4, 16'd55};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 55, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6337] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6338] = {5'd0, 4'd8, 4'd0, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 10, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6339] = {5'd1, 4'd2, 4'd4, 16'd56};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 56, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6340] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6341] = {5'd0, 4'd8, 4'd0, 16'd83};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 83, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6342] = {5'd1, 4'd2, 4'd4, 16'd57};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 57, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6343] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6344] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6345] = {5'd1, 4'd2, 4'd4, 16'd58};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 58, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6346] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6347] = {5'd0, 4'd8, 4'd0, 16'd114};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 114, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6348] = {5'd1, 4'd2, 4'd4, 16'd59};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 59, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6349] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6350] = {5'd0, 4'd8, 4'd0, 16'd118};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 118, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6351] = {5'd1, 4'd2, 4'd4, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 60, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6352] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6353] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6354] = {5'd1, 4'd2, 4'd4, 16'd61};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 61, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6355] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6356] = {5'd0, 4'd8, 4'd0, 16'd114};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 114, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6357] = {5'd1, 4'd2, 4'd4, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 62, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6358] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6359] = {5'd0, 4'd8, 4'd0, 16'd58};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 58, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6360] = {5'd1, 4'd2, 4'd4, 16'd63};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 63, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6361] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6362] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6363] = {5'd1, 4'd2, 4'd4, 16'd64};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 64, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6364] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6365] = {5'd0, 4'd8, 4'd0, 16'd99};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 99, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6366] = {5'd1, 4'd2, 4'd4, 16'd65};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 65, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6367] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6368] = {5'd0, 4'd8, 4'd0, 16'd104};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 104, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6369] = {5'd1, 4'd2, 4'd4, 16'd66};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 66, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6370] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6371] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6372] = {5'd1, 4'd2, 4'd4, 16'd67};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 67, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6373] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6374] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6375] = {5'd1, 4'd2, 4'd4, 16'd68};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 68, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6376] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6377] = {5'd0, 4'd8, 4'd0, 16'd115};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 115, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6378] = {5'd1, 4'd2, 4'd4, 16'd69};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 69, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6379] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6380] = {5'd0, 4'd8, 4'd0, 16'd45};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 45, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6381] = {5'd1, 4'd2, 4'd4, 16'd70};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 70, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6382] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6383] = {5'd0, 4'd8, 4'd0, 16'd119};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 119, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6384] = {5'd1, 4'd2, 4'd4, 16'd71};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 71, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6385] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6386] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6387] = {5'd1, 4'd2, 4'd4, 16'd72};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 72, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6388] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6389] = {5'd0, 4'd8, 4'd0, 16'd98};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 98, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6390] = {5'd1, 4'd2, 4'd4, 16'd73};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 73, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6391] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6392] = {5'd0, 4'd8, 4'd0, 16'd47};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 47, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6393] = {5'd1, 4'd2, 4'd4, 16'd74};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 74, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6394] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6395] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6396] = {5'd1, 4'd2, 4'd4, 16'd75};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 75, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6397] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6398] = {5'd0, 4'd8, 4'd0, 16'd46};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 46, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6399] = {5'd1, 4'd2, 4'd4, 16'd76};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 76, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6400] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6401] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6402] = {5'd1, 4'd2, 4'd4, 16'd77};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 77, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6403] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6404] = {5'd0, 4'd8, 4'd0, 16'd13};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 13, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6405] = {5'd1, 4'd2, 4'd4, 16'd78};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 78, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6406] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6407] = {5'd0, 4'd8, 4'd0, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 10, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6408] = {5'd1, 4'd2, 4'd4, 16'd79};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 79, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6409] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6410] = {5'd0, 4'd8, 4'd0, 16'd67};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 67, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6411] = {5'd1, 4'd2, 4'd4, 16'd80};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 80, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6412] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6413] = {5'd0, 4'd8, 4'd0, 16'd111};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 111, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6414] = {5'd1, 4'd2, 4'd4, 16'd81};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 81, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6415] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6416] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6417] = {5'd1, 4'd2, 4'd4, 16'd82};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 82, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6418] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6419] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6420] = {5'd1, 4'd2, 4'd4, 16'd83};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 83, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6421] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6422] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6423] = {5'd1, 4'd2, 4'd4, 16'd84};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 84, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6424] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6425] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6426] = {5'd1, 4'd2, 4'd4, 16'd85};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 85, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6427] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6428] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6429] = {5'd1, 4'd2, 4'd4, 16'd86};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 86, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6430] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6431] = {5'd0, 4'd8, 4'd0, 16'd45};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 45, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6432] = {5'd1, 4'd2, 4'd4, 16'd87};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 87, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6433] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6434] = {5'd0, 4'd8, 4'd0, 16'd84};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 84, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6435] = {5'd1, 4'd2, 4'd4, 16'd88};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 88, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6436] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6437] = {5'd0, 4'd8, 4'd0, 16'd121};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 121, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6438] = {5'd1, 4'd2, 4'd4, 16'd89};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 89, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6439] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6440] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6441] = {5'd1, 4'd2, 4'd4, 16'd90};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 90, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6442] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6443] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6444] = {5'd1, 4'd2, 4'd4, 16'd91};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 91, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6445] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6446] = {5'd0, 4'd8, 4'd0, 16'd58};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 58, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6447] = {5'd1, 4'd2, 4'd4, 16'd92};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 92, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6448] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6449] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6450] = {5'd1, 4'd2, 4'd4, 16'd93};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 93, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6451] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6452] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6453] = {5'd1, 4'd2, 4'd4, 16'd94};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 94, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6454] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6455] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6456] = {5'd1, 4'd2, 4'd4, 16'd95};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 95, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6457] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6458] = {5'd0, 4'd8, 4'd0, 16'd120};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 120, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6459] = {5'd1, 4'd2, 4'd4, 16'd96};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 96, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6460] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6461] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6462] = {5'd1, 4'd2, 4'd4, 16'd97};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 97, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6463] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6464] = {5'd0, 4'd8, 4'd0, 16'd47};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 47, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6465] = {5'd1, 4'd2, 4'd4, 16'd98};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 98, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6466] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6467] = {5'd0, 4'd8, 4'd0, 16'd104};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 104, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6468] = {5'd1, 4'd2, 4'd4, 16'd99};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 99, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6469] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6470] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6471] = {5'd1, 4'd2, 4'd4, 16'd100};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 100, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6472] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6473] = {5'd0, 4'd8, 4'd0, 16'd109};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 109, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6474] = {5'd1, 4'd2, 4'd4, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 101, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6475] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6476] = {5'd0, 4'd8, 4'd0, 16'd108};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 108, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6477] = {5'd1, 4'd2, 4'd4, 16'd102};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 102, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6478] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6479] = {5'd0, 4'd8, 4'd0, 16'd13};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 13, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6480] = {5'd1, 4'd2, 4'd4, 16'd103};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 103, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6481] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6482] = {5'd0, 4'd8, 4'd0, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 10, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6483] = {5'd1, 4'd2, 4'd4, 16'd104};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 104, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6484] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6485] = {5'd0, 4'd8, 4'd0, 16'd67};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 67, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6486] = {5'd1, 4'd2, 4'd4, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 105, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6487] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6488] = {5'd0, 4'd8, 4'd0, 16'd111};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 111, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6489] = {5'd1, 4'd2, 4'd4, 16'd106};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 106, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6490] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6491] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6492] = {5'd1, 4'd2, 4'd4, 16'd107};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 107, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6493] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6494] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6495] = {5'd1, 4'd2, 4'd4, 16'd108};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 108, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6496] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6497] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6498] = {5'd1, 4'd2, 4'd4, 16'd109};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 109, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6499] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6500] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6501] = {5'd1, 4'd2, 4'd4, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 110, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6502] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6503] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6504] = {5'd1, 4'd2, 4'd4, 16'd111};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 111, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6505] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6506] = {5'd0, 4'd8, 4'd0, 16'd45};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 45, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6507] = {5'd1, 4'd2, 4'd4, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 112, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6508] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6509] = {5'd0, 4'd8, 4'd0, 16'd76};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 76, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6510] = {5'd1, 4'd2, 4'd4, 16'd113};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 113, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6511] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6512] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6513] = {5'd1, 4'd2, 4'd4, 16'd114};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 114, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6514] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6515] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6516] = {5'd1, 4'd2, 4'd4, 16'd115};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 115, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6517] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6518] = {5'd0, 4'd8, 4'd0, 16'd103};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 103, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6519] = {5'd1, 4'd2, 4'd4, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 116, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6520] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6521] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6522] = {5'd1, 4'd2, 4'd4, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 117, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6523] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6524] = {5'd0, 4'd8, 4'd0, 16'd104};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 104, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6525] = {5'd1, 4'd2, 4'd4, 16'd118};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 118, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6526] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6527] = {5'd0, 4'd8, 4'd0, 16'd58};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 58, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6528] = {5'd1, 4'd2, 4'd4, 16'd119};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 119, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6529] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6530] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6531] = {5'd1, 4'd2, 4'd4, 16'd120};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 120, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6532] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6533] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6534] = {5'd1, 4'd2, 4'd4, 16'd121};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 121, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6535] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6536] = {5'd0, 4'd8, 4'd0, 16'd13};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 13, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6537] = {5'd1, 4'd2, 4'd4, 16'd122};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 122, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6538] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6539] = {5'd0, 4'd8, 4'd0, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 10, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6540] = {5'd1, 4'd2, 4'd4, 16'd123};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 123, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6541] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6542] = {5'd0, 4'd8, 4'd0, 16'd13};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 13, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6543] = {5'd1, 4'd2, 4'd4, 16'd124};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 124, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6544] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6545] = {5'd0, 4'd8, 4'd0, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 10, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6546] = {5'd1, 4'd2, 4'd4, 16'd125};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 125, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6547] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6548] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'literal'}
    instructions[6549] = {5'd1, 4'd2, 4'd4, 16'd126};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 4, 'literal': 126, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'addl'}
    instructions[6550] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 92, 'op': 'store'}
    instructions[6551] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 99 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 99, 'op': 'literal'}
    instructions[6552] = {5'd1, 4'd2, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 99 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 99, 'op': 'addl'}
    instructions[6553] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 99 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 99, 'op': 'store'}
    instructions[6554] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100, 'op': 'addl'}
    instructions[6555] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100, 'op': 'store'}
    instructions[6556] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100, 'op': 'addl'}
    instructions[6557] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100, 'op': 'addl'}
    instructions[6558] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100, 'op': 'addl'}
    instructions[6559] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100, 'op': 'load'}
    instructions[6560] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[6561] = {5'd5, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100, 'op': 'load'}
    instructions[6562] = {5'd11, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100, 'op': 'add'}
    instructions[6563] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100, 'op': 'addl'}
    instructions[6564] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100, 'op': 'load'}
    instructions[6565] = {5'd8, 4'd0, 4'd8, 16'd6585};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 101 {'a': 8, 'label': 6585, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 101, 'op': 'jmp_if_false'}
    instructions[6566] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100, 'op': 'addl'}
    instructions[6567] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100, 'op': 'addl'}
    instructions[6568] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100, 'op': 'load'}
    instructions[6569] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100, 'op': 'store'}
    instructions[6570] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100, 'op': 'addl'}
    instructions[6571] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100, 'op': 'literal'}
    instructions[6572] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100, 'op': 'store'}
    instructions[6573] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100, 'op': 'addl'}
    instructions[6574] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100, 'op': 'addl'}
    instructions[6575] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100, 'op': 'addl'}
    instructions[6576] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100, 'op': 'load'}
    instructions[6577] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[6578] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100, 'op': 'load'}
    instructions[6579] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100, 'op': 'add'}
    instructions[6580] = {5'd1, 4'd2, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100, 'op': 'addl'}
    instructions[6581] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100, 'op': 'store'}
    instructions[6582] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[6583] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100, 'op': 'load'}
    instructions[6584] = {5'd12, 4'd0, 4'd0, 16'd6586};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 101 {'label': 6586, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 101, 'op': 'goto'}
    instructions[6585] = {5'd12, 4'd0, 4'd0, 16'd6587};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 101 {'label': 6587, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 101, 'op': 'goto'}
    instructions[6586] = {5'd12, 4'd0, 4'd0, 16'd6554};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100 {'label': 6554, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 100, 'op': 'goto'}
    instructions[6587] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 101 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 101, 'op': 'store'}
    instructions[6588] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 101 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 101, 'op': 'addl'}
    instructions[6589] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 101 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 101, 'op': 'store'}
    instructions[6590] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 101 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 101, 'op': 'addl'}
    instructions[6591] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 101 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 101, 'op': 'addl'}
    instructions[6592] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 101 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 101, 'op': 'addl'}
    instructions[6593] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 101 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 101, 'op': 'load'}
    instructions[6594] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 101 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 101, 'op': 'store'}
    instructions[6595] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 101 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 101, 'op': 'addl'}
    instructions[6596] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 101 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 101, 'op': 'addl'}
    instructions[6597] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 101 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 101, 'op': 'addl'}
    instructions[6598] = {5'd3, 4'd6, 4'd0, 16'd5537};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 101 {'z': 6, 'label': 5537, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 101, 'op': 'call'}
    instructions[6599] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 101 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 101, 'op': 'addl'}
    instructions[6600] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 101 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 101, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[6601] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 101 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 101, 'op': 'load'}
    instructions[6602] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 101 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 101, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[6603] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 101 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 101, 'op': 'load'}
    instructions[6604] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 101 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 101, 'op': 'addl'}
    instructions[6605] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 102 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 102, 'op': 'store'}
    instructions[6606] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 102 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 102, 'op': 'addl'}
    instructions[6607] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 102 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 102, 'op': 'store'}
    instructions[6608] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 102 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 102, 'op': 'addl'}
    instructions[6609] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 102 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 102, 'op': 'addl'}
    instructions[6610] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 102 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 102, 'op': 'store'}
    instructions[6611] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 102 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 102, 'op': 'addl'}
    instructions[6612] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 102 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 102, 'op': 'addl'}
    instructions[6613] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 102 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 102, 'op': 'addl'}
    instructions[6614] = {5'd3, 4'd6, 4'd0, 16'd5553};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 102 {'z': 6, 'label': 5553, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 102, 'op': 'call'}
    instructions[6615] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 102 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 102, 'op': 'addl'}
    instructions[6616] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 102 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 102, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[6617] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 102 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 102, 'op': 'load'}
    instructions[6618] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 102 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 102, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[6619] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 102 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 102, 'op': 'load'}
    instructions[6620] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 102 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 102, 'op': 'addl'}
    instructions[6621] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 103 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 103, 'op': 'store'}
    instructions[6622] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 103 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 103, 'op': 'addl'}
    instructions[6623] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 103 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 103, 'op': 'store'}
    instructions[6624] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 103 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 103, 'op': 'addl'}
    instructions[6625] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 103 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 103, 'op': 'addl'}
    instructions[6626] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 103 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 103, 'op': 'addl'}
    instructions[6627] = {5'd3, 4'd6, 4'd0, 16'd6136};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 103 {'z': 6, 'label': 6136, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 103, 'op': 'call'}
    instructions[6628] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 103 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 103, 'op': 'addl'}
    instructions[6629] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 103 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 103, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[6630] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 103 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 103, 'op': 'load'}
    instructions[6631] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 103 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 103, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[6632] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 103 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 103, 'op': 'load'}
    instructions[6633] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 103 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 103, 'op': 'addl'}
    instructions[6634] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 89 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 89, 'op': 'addl'}
    instructions[6635] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 89 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 89, 'op': 'addl'}
    instructions[6636] = {5'd19, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 89 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/HTTP.h : 89, 'op': 'return'}
  end

  
  always @(posedge clk)
  begin
    load_data <= memory[load_address];
    if(store_enable && state == execute) begin
      memory[store_address] <= store_data;
    end
  end


  //////////////////////////////////////////////////////////////////////////////
  // PIPELINE STAGE 1 -- FETCH INSTRUCTION
  //                                                                            
  
  always @(posedge clk)
  begin
    //implement memory for instructions
    if (state == instruction_fetch || state == operand_fetch || state == execute) begin
      instruction <= instructions[program_counter];
      program_counter_1 <= program_counter;
    end
  end

  assign opcode    = instruction[28:24];
  assign address_z = instruction[23:20];
  assign address_a = instruction[19:16];
  assign address_b = instruction[3:0];
  assign literal   = instruction[15:0];

  //////////////////////////////////////////////////////////////////////////////
  // PIPELINE STAGE 2 -- FETCH OPERANDS
  //                                                                            
  
  always @(posedge clk)
  begin
    if (write_enable) begin
      registers[address_z_3] <= result;
    end
    if (state == operand_fetch || state == execute) begin
      opcode_2 <= opcode;
      literal_2 <= literal;
      address_a_2 <= address_a;
      address_b_2 <= address_b;
      address_z_2 <= address_z;
      program_counter_2 <= program_counter_1;
    end
  end
  assign register_a = registers[address_a_2];
  assign register_b = registers[address_b_2];
  assign operand_a = (address_a_2 == address_z_3 && write_enable)?result:register_a;
  assign operand_b = (address_b_2 == address_z_3 && write_enable)?result:register_b;
  assign store_address = operand_a;
  assign load_address = operand_a;
  assign store_data = operand_b;
  assign store_enable = (opcode_2==2);

  //////////////////////////////////////////////////////////////////////////////
  // PIPELINE STAGE 3 -- EXECUTE
  //                                                                            
  
  always @(posedge clk)
  begin

  write_enable <= 0;
  timer_clock <= timer_clock + 1;
  case(state)

    //instruction_fetch
    instruction_fetch: begin
      program_counter <= program_counter + 1;
      state <= operand_fetch;
    end
    //operand_fetch
    operand_fetch: begin
      program_counter <= program_counter + 1;
      state <= execute;
    end
    //execute
    execute: begin
      program_counter <= program_counter + 1;
      address_z_3 <= address_z_2;
      case(opcode_2)

        //literal
        16'd0:
        begin
          result<=$signed(literal_2);
          write_enable <= 1;
        end

        //addl
        16'd1:
        begin
          result<=operand_a + literal_2;
          write_enable <= 1;
        end

        //store
        16'd2:
        begin
        end

        //call
        16'd3:
        begin
          result <= program_counter_2 + 1;
          write_enable <= 1;
          program_counter <= literal_2;
          state <= instruction_fetch;
        end

        //stop
        16'd4:
        begin
        state <= stop;
        end

        //load
        16'd5:
        begin
          state <= load;
        end

        //read
        16'd6:
        begin
          state <= read;
          read_input <= operand_a;
        end

        //unsigned_greater
        16'd7:
        begin
          result <= $unsigned(operand_a) > $unsigned(operand_b);
          write_enable <= 1;
        end

        //jmp_if_false
        16'd8:
        begin
          if (operand_a == 0) begin
            program_counter <= literal_2;
            state <= instruction_fetch;
          end
        end

        //unsigned_shift_right
        16'd9:
        begin
          if(operand_b < 32) begin
            result <= operand_a >> operand_b;
            carry <= operand_a << (32-operand_b);
          end else begin
            result <= 0;
            carry <= operand_a;
          end
          write_enable <= 1;
        end

        //and
        16'd10:
        begin
          result <= operand_a & operand_b;
          write_enable <= 1;
        end

        //add
        16'd11:
        begin
          long_result = operand_a + operand_b;
          result <= long_result[31:0];
          carry[0] <= long_result[32];
          write_enable <= 1;
        end

        //goto
        16'd12:
        begin
          program_counter <= literal_2;
          state <= instruction_fetch;
        end

        //equal
        16'd13:
        begin
          result <= operand_a == operand_b;
          write_enable <= 1;
        end

        //jmp_if_true
        16'd14:
        begin
          if (operand_a != 0) begin
            program_counter <= literal_2;
            state <= instruction_fetch;
          end
        end

        //not_equal
        16'd15:
        begin
          result <= operand_a != operand_b;
          write_enable <= 1;
        end

        //or
        16'd16:
        begin
          result <= operand_a | operand_b;
          write_enable <= 1;
        end

        //write
        16'd17:
        begin
          state <= write;
          write_output <= operand_a;
          write_value <= operand_b;
        end

        //not
        16'd18:
        begin
          result <= ~operand_a;
          write_enable <= 1;
        end

        //return
        16'd19:
        begin
          program_counter <= operand_a;
          state <= instruction_fetch;
        end

        //unsigned_greater_equal
        16'd20:
        begin
          result <= $unsigned(operand_a) >= $unsigned(operand_b);
          write_enable <= 1;
        end

        //subtract
        16'd21:
        begin
          long_result = operand_a + (~operand_b) + 1;
          result <= long_result[31:0];
          carry[0] <= ~long_result[32];
          write_enable <= 1;
        end

        //shift_left
        16'd22:
        begin
          if(operand_b < 32) begin
            result <= operand_a << operand_b;
            carry <= operand_a >> (32-operand_b);
          end else begin
            result <= 0;
            carry <= operand_a;
          end
          write_enable <= 1;
        end

      endcase

    end

    read:
    begin
      case(read_input)
      0:
      begin
        s_input_socket_ack <= 1;
        if (s_input_socket_ack && input_socket_stb) begin
          result <= input_socket;
          write_enable <= 1;
          s_input_socket_ack <= 0;
          state <= execute;
        end
      end
      3:
      begin
        s_input_rs232_rx_ack <= 1;
        if (s_input_rs232_rx_ack && input_rs232_rx_stb) begin
          result <= input_rs232_rx;
          write_enable <= 1;
          s_input_rs232_rx_ack <= 0;
          state <= execute;
        end
      end
      4:
      begin
        s_input_switches_ack <= 1;
        if (s_input_switches_ack && input_switches_stb) begin
          result <= input_switches;
          write_enable <= 1;
          s_input_switches_ack <= 0;
          state <= execute;
        end
      end
      5:
      begin
        s_input_buttons_ack <= 1;
        if (s_input_buttons_ack && input_buttons_stb) begin
          result <= input_buttons;
          write_enable <= 1;
          s_input_buttons_ack <= 0;
          state <= execute;
        end
      end
      endcase
    end

    write:
    begin
      case(write_output)
      1:
      begin
        s_output_socket_stb <= 1;
        s_output_socket <= write_value;
        if (output_socket_ack && s_output_socket_stb) begin
          s_output_socket_stb <= 0;
          state <= execute;
        end
      end
      2:
      begin
        s_output_rs232_tx_stb <= 1;
        s_output_rs232_tx <= write_value;
        if (output_rs232_tx_ack && s_output_rs232_tx_stb) begin
          s_output_rs232_tx_stb <= 0;
          state <= execute;
        end
      end
      6:
      begin
        s_output_leds_stb <= 1;
        s_output_leds <= write_value;
        if (output_leds_ack && s_output_leds_stb) begin
          s_output_leds_stb <= 0;
          state <= execute;
        end
      end
      endcase
    end

    load:
    begin
        result <= load_data;
        write_enable <= 1;
        state <= execute;
    end

    wait_state:
    begin
      if (timer) begin
        timer <= timer - 1;
      end else begin
        state <= execute;
      end
    end

    stop:
    begin
    end

    endcase

    if (rst == 1'b1) begin
      timer <= 0;
      timer_clock <= 0;
      program_counter <= 0;
      address_z_3 <= 0;
      result <= 0;
      a = 0;
      b = 0;
      z = 0;
      state <= instruction_fetch;
      s_input_socket_ack <= 0;
      s_input_rs232_rx_ack <= 0;
      s_input_switches_ack <= 0;
      s_input_buttons_ack <= 0;
      s_output_socket_stb <= 0;
      s_output_rs232_tx_stb <= 0;
      s_output_leds_stb <= 0;
    end
  end
  assign input_socket_ack = s_input_socket_ack;
  assign input_rs232_rx_ack = s_input_rs232_rx_ack;
  assign input_switches_ack = s_input_switches_ack;
  assign input_buttons_ack = s_input_buttons_ack;
  assign output_socket_stb = s_output_socket_stb;
  assign output_socket = s_output_socket;
  assign output_rs232_tx_stb = s_output_rs232_tx_stb;
  assign output_rs232_tx = s_output_rs232_tx;
  assign output_leds_stb = s_output_leds_stb;
  assign output_leds = s_output_leds;

endmodule
