//name : main_2
//input : input_eth_rx:16
//input : input_socket:16
//output : output_eth_tx:16
//output : output_socket:16
//output : output_rs232_tx:16
//source_file : /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c

///+============================================================================+
///|                                                                            |
///|                     This file was generated by Chips                       |
///|                                                                            |
///|                                  Chips                                     |
///|                                                                            |
///|                      http://github.com/dawsonjon/Chips-2.0                 |
///|                                                                            |
///|                                                             Python powered |
///+============================================================================+
module main_2(input_eth_rx,input_socket,input_eth_rx_stb,input_socket_stb,output_eth_tx_ack,output_socket_ack,output_rs232_tx_ack,clk,rst,output_eth_tx,output_socket,output_rs232_tx,output_eth_tx_stb,output_socket_stb,output_rs232_tx_stb,input_eth_rx_ack,input_socket_ack,exception);
  integer file_count;
  parameter  stop = 3'd0,
  instruction_fetch = 3'd1,
  operand_fetch = 3'd2,
  execute = 3'd3,
  load = 3'd4,
  wait_state = 3'd5,
  read = 3'd6,
  write = 3'd7;
  input [31:0] input_eth_rx;
  input [31:0] input_socket;
  input input_eth_rx_stb;
  input input_socket_stb;
  input output_eth_tx_ack;
  input output_socket_ack;
  input output_rs232_tx_ack;
  input clk;
  input rst;
  output [31:0] output_eth_tx;
  output [31:0] output_socket;
  output [31:0] output_rs232_tx;
  output output_eth_tx_stb;
  output output_socket_stb;
  output output_rs232_tx_stb;
  output input_eth_rx_ack;
  output input_socket_ack;
  reg [31:0] timer;
  reg [63:0] timer_clock;
  reg [15:0] program_counter;
  reg [15:0] program_counter_1;
  reg [15:0] program_counter_2;
  reg [44:0] instruction;
  reg [4:0] opcode_2;
  reg [3:0] a;
  reg [3:0] b;
  reg [3:0] z;
  reg write_enable;
  reg [3:0] address_a_2;
  reg [3:0] address_b_2;
  reg [3:0] address_z_2;
  reg [3:0] address_z_3;
  reg [31:0] load_data;
  reg [31:0] write_output;
  reg [31:0] write_value;
  reg [31:0] read_input;
  reg [15:0] literal_2;
  reg [31:0] a_hi;
  reg [31:0] b_hi;
  reg [31:0] a_lo;
  reg [31:0] b_lo;
  reg [63:0] long_result;
  reg [31:0] result;
  reg [15:0] address;
  reg [31:0] data_out;
  reg [31:0] data_in;
  reg [31:0] carry;
  reg [31:0] s_output_eth_tx_stb;
  reg [31:0] s_output_socket_stb;
  reg [31:0] s_output_rs232_tx_stb;
  reg [31:0] s_output_eth_tx;
  reg [31:0] s_output_socket;
  reg [31:0] s_output_rs232_tx;
  reg [31:0] s_input_eth_rx_ack;
  reg [31:0] s_input_socket_ack;
  reg [7:0] state;
  output reg exception;
  reg [28:0] instructions [5502:0];
  reg [31:0] memory [4096:0];
  reg [31:0] registers [15:0];
  wire [31:0] operand_a;
  wire [31:0] operand_b;
  wire [31:0] register_a;
  wire [31:0] register_b;
  wire [15:0] literal;
  wire [4:0] opcode;
  wire [3:0] address_a;
  wire [3:0] address_b;
  wire [3:0] address_z;
  wire [15:0] load_address;
  wire [15:0] store_address;
  wire [31:0] store_data;
  wire  store_enable;

  //////////////////////////////////////////////////////////////////////////////
  // INSTRUCTION INITIALIZATION                                                 
  //                                                                            
  // Initialise the contents of the instruction memory                          
  //
  // Intruction Set
  // ==============
  // 0 {'literal': True, 'op': 'literal'}
  // 1 {'literal': True, 'op': 'addl'}
  // 2 {'literal': False, 'op': 'store'}
  // 3 {'literal': True, 'op': 'literal_hi'}
  // 4 {'literal': True, 'op': 'call'}
  // 5 {'literal': False, 'op': 'stop'}
  // 6 {'literal': False, 'op': 'load'}
  // 7 {'literal': False, 'op': 'add'}
  // 8 {'literal': True, 'op': 'jmp_if_false'}
  // 9 {'literal': False, 'op': 'subtract'}
  // 10 {'literal': True, 'op': 'goto'}
  // 11 {'literal': False, 'op': 'equal'}
  // 12 {'literal': True, 'op': 'jmp_if_true'}
  // 13 {'literal': False, 'op': 'not_equal'}
  // 14 {'literal': False, 'op': 'ready'}
  // 15 {'literal': False, 'op': 'wait_clocks'}
  // 16 {'literal': False, 'op': 'return'}
  // 17 {'literal': False, 'op': 'or'}
  // 18 {'literal': False, 'op': 'unsigned_shift_right'}
  // 19 {'literal': False, 'op': 'unsigned_greater'}
  // 20 {'literal': False, 'op': 'int_to_long'}
  // 21 {'literal': False, 'op': 'add_with_carry'}
  // 22 {'literal': False, 'op': 'and'}
  // 23 {'literal': False, 'op': 'not'}
  // 24 {'literal': False, 'op': 'unsigned_greater_equal'}
  // 25 {'literal': False, 'op': 'write'}
  // 26 {'literal': False, 'op': 'read'}
  // 27 {'literal': False, 'op': 'shift_right'}
  // 28 {'literal': False, 'op': 'shift_left'}
  // Intructions
  // ===========
  
  initial
  begin
    instructions[0] = {5'd0, 4'd3, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 677 {'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 677, 'op': 'literal'}
    instructions[1] = {5'd0, 4'd4, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 677 {'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 677, 'op': 'literal'}
    instructions[2] = {5'd1, 4'd3, 4'd3, 16'd655};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 677 {'a': 3, 'literal': 655, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 677, 'op': 'addl'}
    instructions[3] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 373 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 373, 'op': 'literal'}
    instructions[4] = {5'd0, 4'd2, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 373 {'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 373, 'op': 'literal'}
    instructions[5] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 373 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 373, 'op': 'store'}
    instructions[6] = {5'd0, 4'd8, 4'd0, 16'd80};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 25 {'literal': 80, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 25, 'op': 'literal'}
    instructions[7] = {5'd0, 4'd2, 4'd0, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 25 {'literal': 4, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 25, 'op': 'literal'}
    instructions[8] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 25 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 25, 'op': 'store'}
    instructions[9] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 370 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 370, 'op': 'literal'}
    instructions[10] = {5'd0, 4'd2, 4'd0, 16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 370 {'literal': 5, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 370, 'op': 'literal'}
    instructions[11] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 370 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 370, 'op': 'store'}
    instructions[12] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155, 'op': 'literal'}
    instructions[13] = {5'd0, 4'd2, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155 {'literal': 6, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155, 'op': 'literal'}
    instructions[14] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155, 'op': 'store'}
    instructions[15] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155, 'op': 'literal'}
    instructions[16] = {5'd0, 4'd2, 4'd0, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155 {'literal': 7, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155, 'op': 'literal'}
    instructions[17] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155, 'op': 'store'}
    instructions[18] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155, 'op': 'literal'}
    instructions[19] = {5'd0, 4'd2, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155 {'literal': 8, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155, 'op': 'literal'}
    instructions[20] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155, 'op': 'store'}
    instructions[21] = {5'd0, 4'd8, 4'd0, 16'd103};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155 {'literal': 103, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155, 'op': 'literal'}
    instructions[22] = {5'd0, 4'd2, 4'd0, 16'd9};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155 {'literal': 9, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155, 'op': 'literal'}
    instructions[23] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155, 'op': 'store'}
    instructions[24] = {5'd0, 4'd8, 4'd0, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155 {'literal': 10, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155, 'op': 'literal'}
    instructions[25] = {5'd0, 4'd2, 4'd0, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155 {'literal': 10, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155, 'op': 'literal'}
    instructions[26] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155, 'op': 'store'}
    instructions[27] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155, 'op': 'literal'}
    instructions[28] = {5'd0, 4'd2, 4'd0, 16'd11};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155 {'literal': 11, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155, 'op': 'literal'}
    instructions[29] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155, 'op': 'store'}
    instructions[30] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 369 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 369, 'op': 'literal'}
    instructions[31] = {5'd0, 4'd2, 4'd0, 16'd12};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 369 {'literal': 12, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 369, 'op': 'literal'}
    instructions[32] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 369 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 369, 'op': 'store'}
    instructions[33] = {5'd0, 4'd8, 4'd0, 16'd257};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 24 {'literal': 257, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 24, 'op': 'literal'}
    instructions[34] = {5'd0, 4'd2, 4'd0, 16'd13};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 24 {'literal': 13, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 24, 'op': 'literal'}
    instructions[35] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 24 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 24, 'op': 'store'}
    instructions[36] = {5'd0, 4'd8, 4'd0, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 34 {'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 34, 'op': 'literal'}
    instructions[37] = {5'd0, 4'd2, 4'd0, 16'd16};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 34 {'literal': 16, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 34, 'op': 'literal'}
    instructions[38] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 34 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 34, 'op': 'store'}
    instructions[39] = {5'd0, 4'd8, 4'd0, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 35 {'literal': 4, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 35, 'op': 'literal'}
    instructions[40] = {5'd0, 4'd2, 4'd0, 16'd20};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 35 {'literal': 20, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 35, 'op': 'literal'}
    instructions[41] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 35 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 35, 'op': 'store'}
    instructions[42] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 371 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 371, 'op': 'literal'}
    instructions[43] = {5'd0, 4'd2, 4'd0, 16'd22};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 371 {'literal': 22, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 371, 'op': 'literal'}
    instructions[44] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 371 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 371, 'op': 'store'}
    instructions[45] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 363 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 363, 'op': 'literal'}
    instructions[46] = {5'd0, 4'd2, 4'd0, 16'd23};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 363 {'literal': 23, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 363, 'op': 'literal'}
    instructions[47] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 363 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 363, 'op': 'store'}
    instructions[48] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 5 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 5, 'op': 'literal'}
    instructions[49] = {5'd0, 4'd2, 4'd0, 16'd24};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 5 {'literal': 24, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 5, 'op': 'literal'}
    instructions[50] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 5 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 5, 'op': 'store'}
    instructions[51] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 385 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 385, 'op': 'literal'}
    instructions[52] = {5'd0, 4'd2, 4'd0, 16'd25};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 385 {'literal': 25, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 385, 'op': 'literal'}
    instructions[53] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 385 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 385, 'op': 'store'}
    instructions[54] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 20 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 20, 'op': 'literal'}
    instructions[55] = {5'd0, 4'd2, 4'd0, 16'd541};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 20 {'literal': 541, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 20, 'op': 'literal'}
    instructions[56] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 20 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 20, 'op': 'store'}
    instructions[57] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 387 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 387, 'op': 'literal'}
    instructions[58] = {5'd0, 4'd2, 4'd0, 16'd542};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 387 {'literal': 542, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 387, 'op': 'literal'}
    instructions[59] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 387 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 387, 'op': 'store'}
    instructions[60] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 32 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 32, 'op': 'literal'}
    instructions[61] = {5'd0, 4'd2, 4'd0, 16'd544};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 32 {'literal': 544, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 32, 'op': 'literal'}
    instructions[62] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 32 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 32, 'op': 'store'}
    instructions[63] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 386 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 386, 'op': 'literal'}
    instructions[64] = {5'd0, 4'd2, 4'd0, 16'd563};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 386 {'literal': 563, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 386, 'op': 'literal'}
    instructions[65] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 386 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 386, 'op': 'store'}
    instructions[66] = {5'd0, 4'd8, 4'd0, 16'd515};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 21 {'literal': 515, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 21, 'op': 'literal'}
    instructions[67] = {5'd0, 4'd2, 4'd0, 16'd580};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 21 {'literal': 580, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 21, 'op': 'literal'}
    instructions[68] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 21 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 21, 'op': 'store'}
    instructions[69] = {5'd0, 4'd8, 4'd0, 16'd1029};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 22 {'literal': 1029, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 22, 'op': 'literal'}
    instructions[70] = {5'd0, 4'd2, 4'd0, 16'd583};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 22 {'literal': 583, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 22, 'op': 'literal'}
    instructions[71] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 22 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 22, 'op': 'store'}
    instructions[72] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 31 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 31, 'op': 'literal'}
    instructions[73] = {5'd0, 4'd2, 4'd0, 16'd585};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 31 {'literal': 585, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 31, 'op': 'literal'}
    instructions[74] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 31 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 31, 'op': 'store'}
    instructions[75] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 382 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 382, 'op': 'literal'}
    instructions[76] = {5'd0, 4'd2, 4'd0, 16'd586};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 382 {'literal': 586, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 382, 'op': 'literal'}
    instructions[77] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 382 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 382, 'op': 'store'}
    instructions[78] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 384 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 384, 'op': 'literal'}
    instructions[79] = {5'd0, 4'd2, 4'd0, 16'd587};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 384 {'literal': 587, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 384, 'op': 'literal'}
    instructions[80] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 384 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 384, 'op': 'store'}
    instructions[81] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 189 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 189, 'op': 'literal'}
    instructions[82] = {5'd0, 4'd2, 4'd0, 16'd588};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 189 {'literal': 588, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 189, 'op': 'literal'}
    instructions[83] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 189 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 189, 'op': 'store'}
    instructions[84] = {5'd0, 4'd8, 4'd0, 16'd49320};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 23 {'literal': 49320, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 23, 'op': 'literal'}
    instructions[85] = {5'd3, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 23 {'a': 8, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 23, 'op': 'literal_hi'}
    instructions[86] = {5'd0, 4'd2, 4'd0, 16'd590};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 23 {'literal': 590, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 23, 'op': 'literal'}
    instructions[87] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 23 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 23, 'op': 'store'}
    instructions[88] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 362 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 362, 'op': 'literal'}
    instructions[89] = {5'd0, 4'd2, 4'd0, 16'd610};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 362 {'literal': 610, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 362, 'op': 'literal'}
    instructions[90] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 362 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 362, 'op': 'store'}
    instructions[91] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 380 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 380, 'op': 'literal'}
    instructions[92] = {5'd0, 4'd2, 4'd0, 16'd627};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 380 {'literal': 627, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 380, 'op': 'literal'}
    instructions[93] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 380 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 380, 'op': 'store'}
    instructions[94] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 377 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 377, 'op': 'literal'}
    instructions[95] = {5'd0, 4'd2, 4'd0, 16'd628};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 377 {'literal': 628, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 377, 'op': 'literal'}
    instructions[96] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 377 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 377, 'op': 'store'}
    instructions[97] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 383 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 383, 'op': 'literal'}
    instructions[98] = {5'd0, 4'd2, 4'd0, 16'd645};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 383 {'literal': 645, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 383, 'op': 'literal'}
    instructions[99] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 383 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 383, 'op': 'store'}
    instructions[100] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 372 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 372, 'op': 'literal'}
    instructions[101] = {5'd0, 4'd2, 4'd0, 16'd649};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 372 {'literal': 649, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 372, 'op': 'literal'}
    instructions[102] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 372 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 372, 'op': 'store'}
    instructions[103] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 374 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 374, 'op': 'literal'}
    instructions[104] = {5'd0, 4'd2, 4'd0, 16'd650};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 374 {'literal': 650, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 374, 'op': 'literal'}
    instructions[105] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 374 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 374, 'op': 'store'}
    instructions[106] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 376 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 376, 'op': 'literal'}
    instructions[107] = {5'd0, 4'd2, 4'd0, 16'd651};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 376 {'literal': 651, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 376, 'op': 'literal'}
    instructions[108] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 376 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 376, 'op': 'store'}
    instructions[109] = {5'd0, 4'd8, 4'd0, 16'd1460};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 367 {'literal': 1460, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 367, 'op': 'literal'}
    instructions[110] = {5'd0, 4'd2, 4'd0, 16'd653};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 367 {'literal': 653, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 367, 'op': 'literal'}
    instructions[111] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 367 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 367, 'op': 'store'}
    instructions[112] = {5'd0, 4'd8, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 33 {'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 33, 'op': 'literal'}
    instructions[113] = {5'd0, 4'd2, 4'd0, 16'd654};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 33 {'literal': 654, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 33, 'op': 'literal'}
    instructions[114] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 33 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.h : 33, 'op': 'store'}
    instructions[115] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 677 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 677, 'op': 'addl'}
    instructions[116] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 677 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 677, 'op': 'addl'}
    instructions[117] = {5'd4, 4'd6, 4'd0, 16'd119};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 677 {'z': 6, 'label': 119, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 677, 'op': 'call'}
    instructions[118] = {5'd5, 4'd0, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 677 {'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 677, 'op': 'stop'}
    instructions[119] = {5'd1, 4'd3, 4'd3, 16'd2063};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 508 {'a': 3, 'literal': 2063, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 508, 'op': 'addl'}
    instructions[120] = {5'd0, 4'd8, 4'd0, 16'd27};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 512 {'literal': 27, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 512, 'op': 'literal'}
    instructions[121] = {5'd1, 4'd2, 4'd4, 16'd2048};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 512 {'a': 4, 'literal': 2048, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 512, 'op': 'addl'}
    instructions[122] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 512 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 512, 'op': 'store'}
    instructions[123] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 514 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 514, 'op': 'literal'}
    instructions[124] = {5'd1, 4'd2, 4'd4, 16'd2049};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 514 {'a': 4, 'literal': 2049, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 514, 'op': 'addl'}
    instructions[125] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 514 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 514, 'op': 'store'}
    instructions[126] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 515 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 515, 'op': 'literal'}
    instructions[127] = {5'd1, 4'd2, 4'd4, 16'd2050};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 515 {'a': 4, 'literal': 2050, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 515, 'op': 'addl'}
    instructions[128] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 515 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 515, 'op': 'store'}
    instructions[129] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 523 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 523, 'op': 'literal'}
    instructions[130] = {5'd1, 4'd2, 4'd4, 16'd2057};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 523 {'a': 4, 'literal': 2057, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 523, 'op': 'addl'}
    instructions[131] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 523 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 523, 'op': 'store'}
    instructions[132] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 524 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 524, 'op': 'literal'}
    instructions[133] = {5'd1, 4'd2, 4'd4, 16'd2058};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 524 {'a': 4, 'literal': 2058, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 524, 'op': 'addl'}
    instructions[134] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 524 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 524, 'op': 'store'}
    instructions[135] = {5'd0, 4'd8, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 525 {'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 525, 'op': 'literal'}
    instructions[136] = {5'd1, 4'd2, 4'd4, 16'd2059};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 525 {'a': 4, 'literal': 2059, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 525, 'op': 'addl'}
    instructions[137] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 525 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 525, 'op': 'store'}
    instructions[138] = {5'd0, 4'd8, 4'd0, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 526 {'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 526, 'op': 'literal'}
    instructions[139] = {5'd1, 4'd2, 4'd4, 16'd2060};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 526 {'a': 4, 'literal': 2060, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 526, 'op': 'addl'}
    instructions[140] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 526 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 526, 'op': 'store'}
    instructions[141] = {5'd0, 4'd8, 4'd0, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 527 {'literal': 4, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 527, 'op': 'literal'}
    instructions[142] = {5'd1, 4'd2, 4'd4, 16'd2061};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 527 {'a': 4, 'literal': 2061, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 527, 'op': 'addl'}
    instructions[143] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 527 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 527, 'op': 'store'}
    instructions[144] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 528 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 528, 'op': 'literal'}
    instructions[145] = {5'd1, 4'd2, 4'd4, 16'd2062};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 528 {'a': 4, 'literal': 2062, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 528, 'op': 'addl'}
    instructions[146] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 528 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 528, 'op': 'store'}
    instructions[147] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 530 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 530, 'op': 'literal'}
    instructions[148] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 530 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 530, 'op': 'store'}
    instructions[149] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 530 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 530, 'op': 'addl'}
    instructions[150] = {5'd0, 4'd8, 4'd0, 16'd608};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 530 {'literal': 608, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 530, 'op': 'literal'}
    instructions[151] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 530 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 530, 'op': 'store'}
    instructions[152] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 530 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 530, 'op': 'addl'}
    instructions[153] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 530 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 530, 'op': 'literal'}
    instructions[154] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 530 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 530, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[155] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 530 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 530, 'op': 'load'}
    instructions[156] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 530 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 530, 'op': 'add'}
    instructions[157] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 530 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 530, 'op': 'addl'}
    instructions[158] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 530 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 530, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[159] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 530 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 530, 'op': 'load'}
    instructions[160] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 530 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 530, 'op': 'store'}
    instructions[161] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 531 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 531, 'op': 'literal'}
    instructions[162] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 531 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 531, 'op': 'store'}
    instructions[163] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 531 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 531, 'op': 'addl'}
    instructions[164] = {5'd0, 4'd8, 4'd0, 16'd608};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 531 {'literal': 608, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 531, 'op': 'literal'}
    instructions[165] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 531 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 531, 'op': 'store'}
    instructions[166] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 531 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 531, 'op': 'addl'}
    instructions[167] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 531 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 531, 'op': 'literal'}
    instructions[168] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 531 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 531, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[169] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 531 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 531, 'op': 'load'}
    instructions[170] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 531 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 531, 'op': 'add'}
    instructions[171] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 531 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 531, 'op': 'addl'}
    instructions[172] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 531 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 531, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[173] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 531 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 531, 'op': 'load'}
    instructions[174] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 531 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 531, 'op': 'store'}
    instructions[175] = {5'd0, 4'd8, 4'd0, 16'd20};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 533 {'literal': 20, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 533, 'op': 'literal'}
    instructions[176] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 533 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 533, 'op': 'addl'}
    instructions[177] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 533 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 533, 'op': 'load'}
    instructions[178] = {5'd0, 4'd2, 4'd0, 16'd24};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 533 {'literal': 24, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 533, 'op': 'literal'}
    instructions[179] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 533 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 533, 'op': 'store'}
    instructions[180] = {5'd1, 4'd8, 4'd4, 16'd2052};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 538 {'a': 4, 'literal': 2052, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 538, 'op': 'addl'}
    instructions[181] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 538 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 538, 'op': 'addl'}
    instructions[182] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 538 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 538, 'op': 'load'}
    instructions[183] = {5'd8, 4'd0, 4'd8, 16'd203};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 538 {'a': 8, 'label': 203, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 538, 'op': 'jmp_if_false'}
    instructions[184] = {5'd1, 4'd8, 4'd4, 16'd2052};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 539 {'a': 4, 'literal': 2052, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 539, 'op': 'addl'}
    instructions[185] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 539 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 539, 'op': 'addl'}
    instructions[186] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 539 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 539, 'op': 'load'}
    instructions[187] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 539 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 539, 'op': 'store'}
    instructions[188] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 539 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 539, 'op': 'addl'}
    instructions[189] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 539 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 539, 'op': 'literal'}
    instructions[190] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 539 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 539, 'op': 'store'}
    instructions[191] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 539 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 539, 'op': 'addl'}
    instructions[192] = {5'd1, 4'd8, 4'd4, 16'd2052};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 539 {'a': 4, 'literal': 2052, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 539, 'op': 'addl'}
    instructions[193] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 539 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 539, 'op': 'addl'}
    instructions[194] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 539 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 539, 'op': 'load'}
    instructions[195] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 539 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 539, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[196] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 539 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 539, 'op': 'load'}
    instructions[197] = {5'd9, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 539 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 539, 'op': 'subtract'}
    instructions[198] = {5'd1, 4'd2, 4'd4, 16'd2052};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 539 {'a': 4, 'literal': 2052, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 539, 'op': 'addl'}
    instructions[199] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 539 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 539, 'op': 'store'}
    instructions[200] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 539 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 539, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[201] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 539 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 539, 'op': 'load'}
    instructions[202] = {5'd10, 4'd0, 4'd0, 16'd240};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 538 {'label': 240, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 538, 'op': 'goto'}
    instructions[203] = {5'd0, 4'd8, 4'd0, 16'd120};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 541 {'literal': 120, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 541, 'op': 'literal'}
    instructions[204] = {5'd1, 4'd2, 4'd4, 16'd2052};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 541 {'a': 4, 'literal': 2052, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 541, 'op': 'addl'}
    instructions[205] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 541 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 541, 'op': 'store'}
    instructions[206] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 542 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 542, 'op': 'literal'}
    instructions[207] = {5'd1, 4'd2, 4'd4, 16'd2062};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 542 {'a': 4, 'literal': 2062, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 542, 'op': 'addl'}
    instructions[208] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 542 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 542, 'op': 'store'}
    instructions[209] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 543 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 543, 'op': 'literal'}
    instructions[210] = {5'd0, 4'd2, 4'd0, 16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 543 {'literal': 5, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 543, 'op': 'literal'}
    instructions[211] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 543 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 543, 'op': 'store'}
    instructions[212] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 544 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 544, 'op': 'literal'}
    instructions[213] = {5'd0, 4'd2, 4'd0, 16'd12};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 544 {'literal': 12, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 544, 'op': 'literal'}
    instructions[214] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 544 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 544, 'op': 'store'}
    instructions[215] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 545 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 545, 'op': 'literal'}
    instructions[216] = {5'd0, 4'd2, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 545 {'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 545, 'op': 'literal'}
    instructions[217] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 545 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 545, 'op': 'store'}
    instructions[218] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 546 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 546, 'op': 'literal'}
    instructions[219] = {5'd0, 4'd2, 4'd0, 16'd22};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 546 {'literal': 22, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 546, 'op': 'literal'}
    instructions[220] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 546 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 546, 'op': 'store'}
    instructions[221] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 547 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 547, 'op': 'store'}
    instructions[222] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 547 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 547, 'op': 'addl'}
    instructions[223] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 547 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 547, 'op': 'store'}
    instructions[224] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 547 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 547, 'op': 'addl'}
    instructions[225] = {5'd1, 4'd8, 4'd4, 16'd1024};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 547 {'a': 4, 'literal': 1024, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 547, 'op': 'addl'}
    instructions[226] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 547 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 547, 'op': 'store'}
    instructions[227] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 547 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 547, 'op': 'addl'}
    instructions[228] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 547 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 547, 'op': 'literal'}
    instructions[229] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 547 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 547, 'op': 'store'}
    instructions[230] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 547 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 547, 'op': 'addl'}
    instructions[231] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 547 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 547, 'op': 'addl'}
    instructions[232] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 547 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 547, 'op': 'addl'}
    instructions[233] = {5'd4, 4'd6, 4'd0, 16'd1040};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 547 {'z': 6, 'label': 1040, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 547, 'op': 'call'}
    instructions[234] = {5'd1, 4'd3, 4'd3, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 547 {'a': 3, 'literal': -2, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 547, 'op': 'addl'}
    instructions[235] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 547 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 547, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[236] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 547 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 547, 'op': 'load'}
    instructions[237] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 547 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 547, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[238] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 547 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 547, 'op': 'load'}
    instructions[239] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 547 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 547, 'op': 'addl'}
    instructions[240] = {5'd1, 4'd8, 4'd4, 16'd2062};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 551 {'a': 4, 'literal': 2062, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 551, 'op': 'addl'}
    instructions[241] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 551 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 551, 'op': 'addl'}
    instructions[242] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 551 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 551, 'op': 'load'}
    instructions[243] = {5'd0, 4'd0, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 551 {'literal': 0, 'z': 0, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 551, 'op': 'literal'}
    instructions[244] = {5'd11, 4'd0, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 551 {'a': 8, 'b': 0, 'z': 0, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 551, 'op': 'equal'}
    instructions[245] = {5'd12, 4'd0, 4'd0, 16'd259};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 551 {'a': 0, 'label': 259, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 551, 'op': 'jmp_if_true'}
    instructions[246] = {5'd0, 4'd0, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 551 {'literal': 1, 'z': 0, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 551, 'op': 'literal'}
    instructions[247] = {5'd11, 4'd0, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 551 {'a': 8, 'b': 0, 'z': 0, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 551, 'op': 'equal'}
    instructions[248] = {5'd12, 4'd0, 4'd0, 16'd272};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 551 {'a': 0, 'label': 272, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 551, 'op': 'jmp_if_true'}
    instructions[249] = {5'd0, 4'd0, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 551 {'literal': 2, 'z': 0, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 551, 'op': 'literal'}
    instructions[250] = {5'd11, 4'd0, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 551 {'a': 8, 'b': 0, 'z': 0, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 551, 'op': 'equal'}
    instructions[251] = {5'd12, 4'd0, 4'd0, 16'd351};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 551 {'a': 0, 'label': 351, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 551, 'op': 'jmp_if_true'}
    instructions[252] = {5'd0, 4'd0, 4'd0, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 551 {'literal': 3, 'z': 0, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 551, 'op': 'literal'}
    instructions[253] = {5'd11, 4'd0, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 551 {'a': 8, 'b': 0, 'z': 0, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 551, 'op': 'equal'}
    instructions[254] = {5'd12, 4'd0, 4'd0, 16'd472};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 551 {'a': 0, 'label': 472, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 551, 'op': 'jmp_if_true'}
    instructions[255] = {5'd0, 4'd0, 4'd0, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 551 {'literal': 4, 'z': 0, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 551, 'op': 'literal'}
    instructions[256] = {5'd11, 4'd0, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 551 {'a': 8, 'b': 0, 'z': 0, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 551, 'op': 'equal'}
    instructions[257] = {5'd12, 4'd0, 4'd0, 16'd494};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 551 {'a': 0, 'label': 494, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 551, 'op': 'jmp_if_true'}
    instructions[258] = {5'd10, 4'd0, 4'd0, 16'd543};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 551 {'label': 543, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 551, 'op': 'goto'}
    instructions[259] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 553 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 553, 'op': 'literal'}
    instructions[260] = {5'd0, 4'd2, 4'd0, 16'd22};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 553 {'literal': 22, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 553, 'op': 'literal'}
    instructions[261] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 553 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 553, 'op': 'store'}
    instructions[262] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 554 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 554, 'op': 'literal'}
    instructions[263] = {5'd0, 4'd2, 4'd0, 16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 554 {'literal': 5, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 554, 'op': 'literal'}
    instructions[264] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 554 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 554, 'op': 'store'}
    instructions[265] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 555 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 555, 'op': 'literal'}
    instructions[266] = {5'd0, 4'd2, 4'd0, 16'd12};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 555 {'literal': 12, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 555, 'op': 'literal'}
    instructions[267] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 555 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 555, 'op': 'store'}
    instructions[268] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 556 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 556, 'op': 'literal'}
    instructions[269] = {5'd0, 4'd2, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 556 {'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 556, 'op': 'literal'}
    instructions[270] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 556 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 556, 'op': 'store'}
    instructions[271] = {5'd10, 4'd0, 4'd0, 16'd543};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 557 {'label': 543, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 557, 'op': 'goto'}
    instructions[272] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 560 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 560, 'op': 'addl'}
    instructions[273] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 560 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 560, 'op': 'store'}
    instructions[274] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 560 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 560, 'op': 'addl'}
    instructions[275] = {5'd0, 4'd8, 4'd0, 16'd13};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 560 {'literal': 13, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 560, 'op': 'literal'}
    instructions[276] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 560 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 560, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[277] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 560 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 560, 'op': 'load'}
    instructions[278] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 560 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 560, 'op': 'add'}
    instructions[279] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 560 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 560, 'op': 'addl'}
    instructions[280] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 560 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 560, 'op': 'load'}
    instructions[281] = {5'd0, 4'd2, 4'd0, 16'd539};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 560 {'literal': 539, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 560, 'op': 'literal'}
    instructions[282] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 560 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 560, 'op': 'store'}
    instructions[283] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 561 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 561, 'op': 'addl'}
    instructions[284] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 561 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 561, 'op': 'store'}
    instructions[285] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 561 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 561, 'op': 'addl'}
    instructions[286] = {5'd0, 4'd8, 4'd0, 16'd14};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 561 {'literal': 14, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 561, 'op': 'literal'}
    instructions[287] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 561 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 561, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[288] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 561 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 561, 'op': 'load'}
    instructions[289] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 561 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 561, 'op': 'add'}
    instructions[290] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 561 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 561, 'op': 'addl'}
    instructions[291] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 561 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 561, 'op': 'load'}
    instructions[292] = {5'd0, 4'd2, 4'd0, 16'd652};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 561 {'literal': 652, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 561, 'op': 'literal'}
    instructions[293] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 561 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 561, 'op': 'store'}
    instructions[294] = {5'd0, 4'd8, 4'd0, 16'd651};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 562 {'literal': 651, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 562, 'op': 'literal'}
    instructions[295] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 562 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 562, 'op': 'addl'}
    instructions[296] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 562 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 562, 'op': 'load'}
    instructions[297] = {5'd0, 4'd2, 4'd0, 16'd23};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 562 {'literal': 23, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 562, 'op': 'literal'}
    instructions[298] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 562 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 562, 'op': 'store'}
    instructions[299] = {5'd0, 4'd8, 4'd0, 16'd80};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 563 {'literal': 80, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 563, 'op': 'literal'}
    instructions[300] = {5'd0, 4'd2, 4'd0, 16'd610};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 563 {'literal': 610, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 563, 'op': 'literal'}
    instructions[301] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 563 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 563, 'op': 'store'}
    instructions[302] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 565 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 565, 'op': 'store'}
    instructions[303] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 565 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 565, 'op': 'addl'}
    instructions[304] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 565 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 565, 'op': 'store'}
    instructions[305] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 565 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 565, 'op': 'addl'}
    instructions[306] = {5'd0, 4'd8, 4'd0, 16'd561};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 565 {'literal': 561, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 565, 'op': 'literal'}
    instructions[307] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 565 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 565, 'op': 'store'}
    instructions[308] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 565 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 565, 'op': 'addl'}
    instructions[309] = {5'd0, 4'd8, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 565 {'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 565, 'op': 'literal'}
    instructions[310] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 565 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 565, 'op': 'store'}
    instructions[311] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 565 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 565, 'op': 'addl'}
    instructions[312] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 565 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 565, 'op': 'literal'}
    instructions[313] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 565 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 565, 'op': 'store'}
    instructions[314] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 565 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 565, 'op': 'addl'}
    instructions[315] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 565 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 565, 'op': 'addl'}
    instructions[316] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 565 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 565, 'op': 'addl'}
    instructions[317] = {5'd4, 4'd6, 4'd0, 16'd3325};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 565 {'z': 6, 'label': 3325, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 565, 'op': 'call'}
    instructions[318] = {5'd1, 4'd3, 4'd3, -16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 565 {'a': 3, 'literal': -3, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 565, 'op': 'addl'}
    instructions[319] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 565 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 565, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[320] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 565 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 565, 'op': 'load'}
    instructions[321] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 565 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 565, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[322] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 565 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 565, 'op': 'load'}
    instructions[323] = {5'd0, 4'd2, 4'd0, 16'd582};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 565 {'literal': 582, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 565, 'op': 'literal'}
    instructions[324] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 565 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 565, 'op': 'load'}
    instructions[325] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 566 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 566, 'op': 'literal'}
    instructions[326] = {5'd0, 4'd2, 4'd0, 16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 566 {'literal': 5, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 566, 'op': 'literal'}
    instructions[327] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 566 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 566, 'op': 'store'}
    instructions[328] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 567 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 567, 'op': 'literal'}
    instructions[329] = {5'd0, 4'd2, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 567 {'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 567, 'op': 'literal'}
    instructions[330] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 567 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 567, 'op': 'store'}
    instructions[331] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 568 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 568, 'op': 'store'}
    instructions[332] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 568 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 568, 'op': 'addl'}
    instructions[333] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 568 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 568, 'op': 'store'}
    instructions[334] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 568 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 568, 'op': 'addl'}
    instructions[335] = {5'd1, 4'd8, 4'd4, 16'd1024};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 568 {'a': 4, 'literal': 1024, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 568, 'op': 'addl'}
    instructions[336] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 568 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 568, 'op': 'store'}
    instructions[337] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 568 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 568, 'op': 'addl'}
    instructions[338] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 568 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 568, 'op': 'literal'}
    instructions[339] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 568 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 568, 'op': 'store'}
    instructions[340] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 568 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 568, 'op': 'addl'}
    instructions[341] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 568 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 568, 'op': 'addl'}
    instructions[342] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 568 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 568, 'op': 'addl'}
    instructions[343] = {5'd4, 4'd6, 4'd0, 16'd1040};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 568 {'z': 6, 'label': 1040, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 568, 'op': 'call'}
    instructions[344] = {5'd1, 4'd3, 4'd3, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 568 {'a': 3, 'literal': -2, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 568, 'op': 'addl'}
    instructions[345] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 568 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 568, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[346] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 568 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 568, 'op': 'load'}
    instructions[347] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 568 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 568, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[348] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 568 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 568, 'op': 'load'}
    instructions[349] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 568 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 568, 'op': 'addl'}
    instructions[350] = {5'd10, 4'd0, 4'd0, 16'd543};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 569 {'label': 543, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 569, 'op': 'goto'}
    instructions[351] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572, 'op': 'store'}
    instructions[352] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572, 'op': 'addl'}
    instructions[353] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572, 'op': 'store'}
    instructions[354] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572, 'op': 'addl'}
    instructions[355] = {5'd1, 4'd8, 4'd4, 16'd1024};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572 {'a': 4, 'literal': 1024, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572, 'op': 'addl'}
    instructions[356] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572, 'op': 'store'}
    instructions[357] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572, 'op': 'addl'}
    instructions[358] = {5'd1, 4'd8, 4'd4, 16'd2048};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572 {'a': 4, 'literal': 2048, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572, 'op': 'addl'}
    instructions[359] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572, 'op': 'addl'}
    instructions[360] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572, 'op': 'load'}
    instructions[361] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572, 'op': 'store'}
    instructions[362] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572, 'op': 'addl'}
    instructions[363] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572, 'op': 'addl'}
    instructions[364] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572, 'op': 'addl'}
    instructions[365] = {5'd4, 4'd6, 4'd0, 16'd3474};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572 {'z': 6, 'label': 3474, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572, 'op': 'call'}
    instructions[366] = {5'd1, 4'd3, 4'd3, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572 {'a': 3, 'literal': -2, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572, 'op': 'addl'}
    instructions[367] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[368] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572, 'op': 'load'}
    instructions[369] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[370] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572, 'op': 'load'}
    instructions[371] = {5'd0, 4'd2, 4'd0, 16'd543};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572 {'literal': 543, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572, 'op': 'literal'}
    instructions[372] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572, 'op': 'load'}
    instructions[373] = {5'd1, 4'd2, 4'd4, 16'd2051};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572 {'a': 4, 'literal': 2051, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572, 'op': 'addl'}
    instructions[374] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 572, 'op': 'store'}
    instructions[375] = {5'd0, 4'd8, 4'd0, 16'd14};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 573 {'literal': 14, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 573, 'op': 'literal'}
    instructions[376] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 573 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 573, 'op': 'store'}
    instructions[377] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 573 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 573, 'op': 'addl'}
    instructions[378] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 573 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 573, 'op': 'literal'}
    instructions[379] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 573 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 573, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[380] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 573 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 573, 'op': 'load'}
    instructions[381] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 573 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 573, 'op': 'add'}
    instructions[382] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 573 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 573, 'op': 'addl'}
    instructions[383] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 573 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 573, 'op': 'load'}
    instructions[384] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 573 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 573, 'op': 'store'}
    instructions[385] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 573 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 573, 'op': 'addl'}
    instructions[386] = {5'd0, 4'd8, 4'd0, 16'd608};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 573 {'literal': 608, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 573, 'op': 'literal'}
    instructions[387] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 573 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 573, 'op': 'store'}
    instructions[388] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 573 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 573, 'op': 'addl'}
    instructions[389] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 573 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 573, 'op': 'literal'}
    instructions[390] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 573 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 573, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[391] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 573 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 573, 'op': 'load'}
    instructions[392] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 573 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 573, 'op': 'add'}
    instructions[393] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 573 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 573, 'op': 'addl'}
    instructions[394] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 573 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 573, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[395] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 573 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 573, 'op': 'load'}
    instructions[396] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 573 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 573, 'op': 'store'}
    instructions[397] = {5'd0, 4'd8, 4'd0, 16'd14};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 574 {'literal': 14, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 574, 'op': 'literal'}
    instructions[398] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 574 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 574, 'op': 'store'}
    instructions[399] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 574 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 574, 'op': 'addl'}
    instructions[400] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 574 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 574, 'op': 'literal'}
    instructions[401] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 574 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 574, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[402] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 574 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 574, 'op': 'load'}
    instructions[403] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 574 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 574, 'op': 'add'}
    instructions[404] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 574 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 574, 'op': 'addl'}
    instructions[405] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 574 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 574, 'op': 'load'}
    instructions[406] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 574 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 574, 'op': 'store'}
    instructions[407] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 574 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 574, 'op': 'addl'}
    instructions[408] = {5'd0, 4'd8, 4'd0, 16'd608};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 574 {'literal': 608, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 574, 'op': 'literal'}
    instructions[409] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 574 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 574, 'op': 'store'}
    instructions[410] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 574 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 574, 'op': 'addl'}
    instructions[411] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 574 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 574, 'op': 'literal'}
    instructions[412] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 574 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 574, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[413] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 574 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 574, 'op': 'load'}
    instructions[414] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 574 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 574, 'op': 'add'}
    instructions[415] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 574 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 574, 'op': 'addl'}
    instructions[416] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 574 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 574, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[417] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 574 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 574, 'op': 'load'}
    instructions[418] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 574 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 574, 'op': 'store'}
    instructions[419] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575, 'op': 'store'}
    instructions[420] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575, 'op': 'addl'}
    instructions[421] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575, 'op': 'store'}
    instructions[422] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575, 'op': 'addl'}
    instructions[423] = {5'd0, 4'd8, 4'd0, 16'd14};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575 {'literal': 14, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575, 'op': 'literal'}
    instructions[424] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575, 'op': 'store'}
    instructions[425] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575, 'op': 'addl'}
    instructions[426] = {5'd0, 4'd8, 4'd0, 16'd608};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575 {'literal': 608, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575, 'op': 'literal'}
    instructions[427] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575, 'op': 'store'}
    instructions[428] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575, 'op': 'addl'}
    instructions[429] = {5'd1, 4'd8, 4'd4, 16'd2051};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575 {'a': 4, 'literal': 2051, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575, 'op': 'addl'}
    instructions[430] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575, 'op': 'addl'}
    instructions[431] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575, 'op': 'load'}
    instructions[432] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575, 'op': 'store'}
    instructions[433] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575, 'op': 'addl'}
    instructions[434] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575, 'op': 'addl'}
    instructions[435] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575, 'op': 'addl'}
    instructions[436] = {5'd4, 4'd6, 4'd0, 16'd3325};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575 {'z': 6, 'label': 3325, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575, 'op': 'call'}
    instructions[437] = {5'd1, 4'd3, 4'd3, -16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575 {'a': 3, 'literal': -3, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575, 'op': 'addl'}
    instructions[438] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[439] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575, 'op': 'load'}
    instructions[440] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[441] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575, 'op': 'load'}
    instructions[442] = {5'd0, 4'd2, 4'd0, 16'd582};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575 {'literal': 582, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575, 'op': 'literal'}
    instructions[443] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 575, 'op': 'load'}
    instructions[444] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 576 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 576, 'op': 'literal'}
    instructions[445] = {5'd0, 4'd2, 4'd0, 16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 576 {'literal': 5, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 576, 'op': 'literal'}
    instructions[446] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 576 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 576, 'op': 'store'}
    instructions[447] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 577 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 577, 'op': 'literal'}
    instructions[448] = {5'd0, 4'd2, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 577 {'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 577, 'op': 'literal'}
    instructions[449] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 577 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 577, 'op': 'store'}
    instructions[450] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 578 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 578, 'op': 'store'}
    instructions[451] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 578 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 578, 'op': 'addl'}
    instructions[452] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 578 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 578, 'op': 'store'}
    instructions[453] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 578 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 578, 'op': 'addl'}
    instructions[454] = {5'd1, 4'd8, 4'd4, 16'd1024};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 578 {'a': 4, 'literal': 1024, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 578, 'op': 'addl'}
    instructions[455] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 578 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 578, 'op': 'store'}
    instructions[456] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 578 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 578, 'op': 'addl'}
    instructions[457] = {5'd1, 4'd8, 4'd4, 16'd2051};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 578 {'a': 4, 'literal': 2051, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 578, 'op': 'addl'}
    instructions[458] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 578 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 578, 'op': 'addl'}
    instructions[459] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 578 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 578, 'op': 'load'}
    instructions[460] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 578 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 578, 'op': 'store'}
    instructions[461] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 578 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 578, 'op': 'addl'}
    instructions[462] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 578 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 578, 'op': 'addl'}
    instructions[463] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 578 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 578, 'op': 'addl'}
    instructions[464] = {5'd4, 4'd6, 4'd0, 16'd1040};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 578 {'z': 6, 'label': 1040, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 578, 'op': 'call'}
    instructions[465] = {5'd1, 4'd3, 4'd3, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 578 {'a': 3, 'literal': -2, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 578, 'op': 'addl'}
    instructions[466] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 578 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 578, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[467] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 578 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 578, 'op': 'load'}
    instructions[468] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 578 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 578, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[469] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 578 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 578, 'op': 'load'}
    instructions[470] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 578 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 578, 'op': 'addl'}
    instructions[471] = {5'd10, 4'd0, 4'd0, 16'd543};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 579 {'label': 543, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 579, 'op': 'goto'}
    instructions[472] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 582 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 582, 'op': 'store'}
    instructions[473] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 582 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 582, 'op': 'addl'}
    instructions[474] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 582 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 582, 'op': 'store'}
    instructions[475] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 582 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 582, 'op': 'addl'}
    instructions[476] = {5'd1, 4'd8, 4'd4, 16'd1024};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 582 {'a': 4, 'literal': 1024, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 582, 'op': 'addl'}
    instructions[477] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 582 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 582, 'op': 'store'}
    instructions[478] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 582 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 582, 'op': 'addl'}
    instructions[479] = {5'd1, 4'd8, 4'd4, 16'd2051};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 582 {'a': 4, 'literal': 2051, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 582, 'op': 'addl'}
    instructions[480] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 582 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 582, 'op': 'addl'}
    instructions[481] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 582 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 582, 'op': 'load'}
    instructions[482] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 582 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 582, 'op': 'store'}
    instructions[483] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 582 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 582, 'op': 'addl'}
    instructions[484] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 582 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 582, 'op': 'addl'}
    instructions[485] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 582 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 582, 'op': 'addl'}
    instructions[486] = {5'd4, 4'd6, 4'd0, 16'd1040};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 582 {'z': 6, 'label': 1040, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 582, 'op': 'call'}
    instructions[487] = {5'd1, 4'd3, 4'd3, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 582 {'a': 3, 'literal': -2, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 582, 'op': 'addl'}
    instructions[488] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 582 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 582, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[489] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 582 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 582, 'op': 'load'}
    instructions[490] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 582 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 582, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[491] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 582 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 582, 'op': 'load'}
    instructions[492] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 582 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 582, 'op': 'addl'}
    instructions[493] = {5'd10, 4'd0, 4'd0, 16'd543};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 583 {'label': 543, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 583, 'op': 'goto'}
    instructions[494] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 586 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 586, 'op': 'literal'}
    instructions[495] = {5'd0, 4'd2, 4'd0, 16'd12};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 586 {'literal': 12, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 586, 'op': 'literal'}
    instructions[496] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 586 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 586, 'op': 'store'}
    instructions[497] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 587 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 587, 'op': 'literal'}
    instructions[498] = {5'd0, 4'd2, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 587 {'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 587, 'op': 'literal'}
    instructions[499] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 587 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 587, 'op': 'store'}
    instructions[500] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 588 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 588, 'op': 'store'}
    instructions[501] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 588 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 588, 'op': 'addl'}
    instructions[502] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 588 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 588, 'op': 'store'}
    instructions[503] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 588 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 588, 'op': 'addl'}
    instructions[504] = {5'd0, 4'd8, 4'd0, 16'd561};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 588 {'literal': 561, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 588, 'op': 'literal'}
    instructions[505] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 588 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 588, 'op': 'store'}
    instructions[506] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 588 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 588, 'op': 'addl'}
    instructions[507] = {5'd0, 4'd8, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 588 {'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 588, 'op': 'literal'}
    instructions[508] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 588 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 588, 'op': 'store'}
    instructions[509] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 588 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 588, 'op': 'addl'}
    instructions[510] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 588 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 588, 'op': 'literal'}
    instructions[511] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 588 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 588, 'op': 'store'}
    instructions[512] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 588 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 588, 'op': 'addl'}
    instructions[513] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 588 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 588, 'op': 'addl'}
    instructions[514] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 588 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 588, 'op': 'addl'}
    instructions[515] = {5'd4, 4'd6, 4'd0, 16'd3325};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 588 {'z': 6, 'label': 3325, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 588, 'op': 'call'}
    instructions[516] = {5'd1, 4'd3, 4'd3, -16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 588 {'a': 3, 'literal': -3, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 588, 'op': 'addl'}
    instructions[517] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 588 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 588, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[518] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 588 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 588, 'op': 'load'}
    instructions[519] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 588 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 588, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[520] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 588 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 588, 'op': 'load'}
    instructions[521] = {5'd0, 4'd2, 4'd0, 16'd582};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 588 {'literal': 582, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 588, 'op': 'literal'}
    instructions[522] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 588 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 588, 'op': 'load'}
    instructions[523] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 589 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 589, 'op': 'store'}
    instructions[524] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 589 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 589, 'op': 'addl'}
    instructions[525] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 589 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 589, 'op': 'store'}
    instructions[526] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 589 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 589, 'op': 'addl'}
    instructions[527] = {5'd1, 4'd8, 4'd4, 16'd1024};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 589 {'a': 4, 'literal': 1024, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 589, 'op': 'addl'}
    instructions[528] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 589 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 589, 'op': 'store'}
    instructions[529] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 589 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 589, 'op': 'addl'}
    instructions[530] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 589 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 589, 'op': 'literal'}
    instructions[531] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 589 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 589, 'op': 'store'}
    instructions[532] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 589 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 589, 'op': 'addl'}
    instructions[533] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 589 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 589, 'op': 'addl'}
    instructions[534] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 589 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 589, 'op': 'addl'}
    instructions[535] = {5'd4, 4'd6, 4'd0, 16'd1040};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 589 {'z': 6, 'label': 1040, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 589, 'op': 'call'}
    instructions[536] = {5'd1, 4'd3, 4'd3, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 589 {'a': 3, 'literal': -2, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 589, 'op': 'addl'}
    instructions[537] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 589 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 589, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[538] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 589 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 589, 'op': 'load'}
    instructions[539] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 589 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 589, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[540] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 589 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 589, 'op': 'load'}
    instructions[541] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 589 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 589, 'op': 'addl'}
    instructions[542] = {5'd10, 4'd0, 4'd0, 16'd543};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 590 {'label': 543, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 590, 'op': 'goto'}
    instructions[543] = {5'd0, 4'd8, 4'd0, 16'd10000};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594 {'literal': 10000, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594, 'op': 'literal'}
    instructions[544] = {5'd1, 4'd2, 4'd4, 16'd2053};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594 {'a': 4, 'literal': 2053, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594, 'op': 'addl'}
    instructions[545] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594, 'op': 'store'}
    instructions[546] = {5'd1, 4'd8, 4'd4, 16'd2053};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594 {'a': 4, 'literal': 2053, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594, 'op': 'addl'}
    instructions[547] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594, 'op': 'addl'}
    instructions[548] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594, 'op': 'load'}
    instructions[549] = {5'd8, 4'd0, 4'd8, 16'd1036};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594 {'a': 8, 'label': 1036, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594, 'op': 'jmp_if_false'}
    instructions[550] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 595 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 595, 'op': 'store'}
    instructions[551] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 595 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 595, 'op': 'addl'}
    instructions[552] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 595 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 595, 'op': 'store'}
    instructions[553] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 595 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 595, 'op': 'addl'}
    instructions[554] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 595 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 595, 'op': 'addl'}
    instructions[555] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 595 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 595, 'op': 'store'}
    instructions[556] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 595 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 595, 'op': 'addl'}
    instructions[557] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 595 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 595, 'op': 'addl'}
    instructions[558] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 595 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 595, 'op': 'addl'}
    instructions[559] = {5'd4, 4'd6, 4'd0, 16'd3608};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 595 {'z': 6, 'label': 3608, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 595, 'op': 'call'}
    instructions[560] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 595 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 595, 'op': 'addl'}
    instructions[561] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 595 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 595, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[562] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 595 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 595, 'op': 'load'}
    instructions[563] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 595 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 595, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[564] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 595 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 595, 'op': 'load'}
    instructions[565] = {5'd0, 4'd2, 4'd0, 16'd646};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 595 {'literal': 646, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 595, 'op': 'literal'}
    instructions[566] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 595 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 595, 'op': 'load'}
    instructions[567] = {5'd1, 4'd2, 4'd4, 16'd2054};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 595 {'a': 4, 'literal': 2054, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 595, 'op': 'addl'}
    instructions[568] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 595 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 595, 'op': 'store'}
    instructions[569] = {5'd1, 4'd8, 4'd4, 16'd2054};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 596 {'a': 4, 'literal': 2054, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 596, 'op': 'addl'}
    instructions[570] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 596 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 596, 'op': 'addl'}
    instructions[571] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 596 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 596, 'op': 'load'}
    instructions[572] = {5'd8, 4'd0, 4'd8, 16'd582};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 596 {'a': 8, 'label': 582, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 596, 'op': 'jmp_if_false'}
    instructions[573] = {5'd0, 4'd8, 4'd0, 16'd80};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 596 {'literal': 80, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 596, 'op': 'literal'}
    instructions[574] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 596 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 596, 'op': 'store'}
    instructions[575] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 596 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 596, 'op': 'addl'}
    instructions[576] = {5'd0, 4'd8, 4'd0, 16'd628};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 596 {'literal': 628, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 596, 'op': 'literal'}
    instructions[577] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 596 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 596, 'op': 'addl'}
    instructions[578] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 596 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 596, 'op': 'load'}
    instructions[579] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 596 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 596, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[580] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 596 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 596, 'op': 'load'}
    instructions[581] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 596 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 596, 'op': 'equal'}
    instructions[582] = {5'd8, 4'd0, 4'd8, 16'd1015};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 596 {'a': 8, 'label': 1015, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 596, 'op': 'jmp_if_false'}
    instructions[583] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598, 'op': 'literal'}
    instructions[584] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598, 'op': 'store'}
    instructions[585] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598, 'op': 'addl'}
    instructions[586] = {5'd1, 4'd8, 4'd4, 16'd2062};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598 {'a': 4, 'literal': 2062, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598, 'op': 'addl'}
    instructions[587] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598, 'op': 'addl'}
    instructions[588] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598, 'op': 'load'}
    instructions[589] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[590] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598, 'op': 'load'}
    instructions[591] = {5'd13, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598, 'op': 'not_equal'}
    instructions[592] = {5'd8, 4'd0, 4'd8, 16'd604};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598 {'a': 8, 'label': 604, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598, 'op': 'jmp_if_false'}
    instructions[593] = {5'd0, 4'd8, 4'd0, 16'd23};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598 {'literal': 23, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598, 'op': 'literal'}
    instructions[594] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598, 'op': 'addl'}
    instructions[595] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598, 'op': 'load'}
    instructions[596] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598, 'op': 'store'}
    instructions[597] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598, 'op': 'addl'}
    instructions[598] = {5'd0, 4'd8, 4'd0, 16'd651};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598 {'literal': 651, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598, 'op': 'literal'}
    instructions[599] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598, 'op': 'addl'}
    instructions[600] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598, 'op': 'load'}
    instructions[601] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[602] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598, 'op': 'load'}
    instructions[603] = {5'd13, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598, 'op': 'not_equal'}
    instructions[604] = {5'd8, 4'd0, 4'd8, 16'd607};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598 {'a': 8, 'label': 607, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598, 'op': 'jmp_if_false'}
    instructions[605] = {5'd10, 4'd0, 4'd0, 16'd1017};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598 {'label': 1017, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598, 'op': 'goto'}
    instructions[606] = {5'd10, 4'd0, 4'd0, 16'd607};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598 {'label': 607, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 598, 'op': 'goto'}
    instructions[607] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 599 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 599, 'op': 'literal'}
    instructions[608] = {5'd1, 4'd2, 4'd4, 16'd2056};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 599 {'a': 4, 'literal': 2056, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 599, 'op': 'addl'}
    instructions[609] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 599 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 599, 'op': 'store'}
    instructions[610] = {5'd1, 4'd8, 4'd4, 16'd2062};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 600 {'a': 4, 'literal': 2062, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 600, 'op': 'addl'}
    instructions[611] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 600 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 600, 'op': 'addl'}
    instructions[612] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 600 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 600, 'op': 'load'}
    instructions[613] = {5'd1, 4'd2, 4'd4, 16'd2055};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 600 {'a': 4, 'literal': 2055, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 600, 'op': 'addl'}
    instructions[614] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 600 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 600, 'op': 'store'}
    instructions[615] = {5'd1, 4'd8, 4'd4, 16'd2062};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 601 {'a': 4, 'literal': 2062, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 601, 'op': 'addl'}
    instructions[616] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 601 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 601, 'op': 'addl'}
    instructions[617] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 601 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 601, 'op': 'load'}
    instructions[618] = {5'd0, 4'd0, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 601 {'literal': 0, 'z': 0, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 601, 'op': 'literal'}
    instructions[619] = {5'd11, 4'd0, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 601 {'a': 8, 'b': 0, 'z': 0, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 601, 'op': 'equal'}
    instructions[620] = {5'd12, 4'd0, 4'd0, 16'd634};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 601 {'a': 0, 'label': 634, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 601, 'op': 'jmp_if_true'}
    instructions[621] = {5'd0, 4'd0, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 601 {'literal': 1, 'z': 0, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 601, 'op': 'literal'}
    instructions[622] = {5'd11, 4'd0, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 601 {'a': 8, 'b': 0, 'z': 0, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 601, 'op': 'equal'}
    instructions[623] = {5'd12, 4'd0, 4'd0, 16'd665};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 601 {'a': 0, 'label': 665, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 601, 'op': 'jmp_if_true'}
    instructions[624] = {5'd0, 4'd0, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 601 {'literal': 2, 'z': 0, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 601, 'op': 'literal'}
    instructions[625] = {5'd11, 4'd0, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 601 {'a': 8, 'b': 0, 'z': 0, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 601, 'op': 'equal'}
    instructions[626] = {5'd12, 4'd0, 4'd0, 16'd762};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 601 {'a': 0, 'label': 762, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 601, 'op': 'jmp_if_true'}
    instructions[627] = {5'd0, 4'd0, 4'd0, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 601 {'literal': 3, 'z': 0, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 601, 'op': 'literal'}
    instructions[628] = {5'd11, 4'd0, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 601 {'a': 8, 'b': 0, 'z': 0, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 601, 'op': 'equal'}
    instructions[629] = {5'd12, 4'd0, 4'd0, 16'd806};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 601 {'a': 0, 'label': 806, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 601, 'op': 'jmp_if_true'}
    instructions[630] = {5'd0, 4'd0, 4'd0, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 601 {'literal': 4, 'z': 0, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 601, 'op': 'literal'}
    instructions[631] = {5'd11, 4'd0, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 601 {'a': 8, 'b': 0, 'z': 0, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 601, 'op': 'equal'}
    instructions[632] = {5'd12, 4'd0, 4'd0, 16'd898};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 601 {'a': 0, 'label': 898, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 601, 'op': 'jmp_if_true'}
    instructions[633] = {5'd10, 4'd0, 4'd0, 16'd907};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 601 {'label': 907, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 601, 'op': 'goto'}
    instructions[634] = {5'd0, 4'd8, 4'd0, 16'd645};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 605 {'literal': 645, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 605, 'op': 'literal'}
    instructions[635] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 605 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 605, 'op': 'addl'}
    instructions[636] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 605 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 605, 'op': 'load'}
    instructions[637] = {5'd8, 4'd0, 4'd8, 16'd642};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 605 {'a': 8, 'label': 642, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 605, 'op': 'jmp_if_false'}
    instructions[638] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 605 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 605, 'op': 'literal'}
    instructions[639] = {5'd1, 4'd2, 4'd4, 16'd2062};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 605 {'a': 4, 'literal': 2062, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 605, 'op': 'addl'}
    instructions[640] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 605 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 605, 'op': 'store'}
    instructions[641] = {5'd10, 4'd0, 4'd0, 16'd664};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 605 {'label': 664, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 605, 'op': 'goto'}
    instructions[642] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 607 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 607, 'op': 'literal'}
    instructions[643] = {5'd0, 4'd2, 4'd0, 16'd22};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 607 {'literal': 22, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 607, 'op': 'literal'}
    instructions[644] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 607 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 607, 'op': 'store'}
    instructions[645] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 608 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 608, 'op': 'store'}
    instructions[646] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 608 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 608, 'op': 'addl'}
    instructions[647] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 608 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 608, 'op': 'store'}
    instructions[648] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 608 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 608, 'op': 'addl'}
    instructions[649] = {5'd1, 4'd8, 4'd4, 16'd1024};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 608 {'a': 4, 'literal': 1024, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 608, 'op': 'addl'}
    instructions[650] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 608 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 608, 'op': 'store'}
    instructions[651] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 608 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 608, 'op': 'addl'}
    instructions[652] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 608 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 608, 'op': 'literal'}
    instructions[653] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 608 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 608, 'op': 'store'}
    instructions[654] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 608 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 608, 'op': 'addl'}
    instructions[655] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 608 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 608, 'op': 'addl'}
    instructions[656] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 608 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 608, 'op': 'addl'}
    instructions[657] = {5'd4, 4'd6, 4'd0, 16'd1040};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 608 {'z': 6, 'label': 1040, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 608, 'op': 'call'}
    instructions[658] = {5'd1, 4'd3, 4'd3, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 608 {'a': 3, 'literal': -2, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 608, 'op': 'addl'}
    instructions[659] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 608 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 608, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[660] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 608 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 608, 'op': 'load'}
    instructions[661] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 608 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 608, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[662] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 608 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 608, 'op': 'load'}
    instructions[663] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 608 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 608, 'op': 'addl'}
    instructions[664] = {5'd10, 4'd0, 4'd0, 16'd907};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 610 {'label': 907, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 610, 'op': 'goto'}
    instructions[665] = {5'd0, 4'd8, 4'd0, 16'd563};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 614 {'literal': 563, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 614, 'op': 'literal'}
    instructions[666] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 614 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 614, 'op': 'addl'}
    instructions[667] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 614 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 614, 'op': 'load'}
    instructions[668] = {5'd8, 4'd0, 4'd8, 16'd761};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 614 {'a': 8, 'label': 761, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 614, 'op': 'jmp_if_false'}
    instructions[669] = {5'd0, 4'd8, 4'd0, 16'd18};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 615 {'literal': 18, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 615, 'op': 'literal'}
    instructions[670] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 615 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 615, 'op': 'store'}
    instructions[671] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 615 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 615, 'op': 'addl'}
    instructions[672] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 615 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 615, 'op': 'literal'}
    instructions[673] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 615 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 615, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[674] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 615 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 615, 'op': 'load'}
    instructions[675] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 615 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 615, 'op': 'add'}
    instructions[676] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 615 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 615, 'op': 'addl'}
    instructions[677] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 615 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 615, 'op': 'load'}
    instructions[678] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 615 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 615, 'op': 'store'}
    instructions[679] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 615 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 615, 'op': 'addl'}
    instructions[680] = {5'd0, 4'd8, 4'd0, 16'd608};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 615 {'literal': 608, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 615, 'op': 'literal'}
    instructions[681] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 615 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 615, 'op': 'store'}
    instructions[682] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 615 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 615, 'op': 'addl'}
    instructions[683] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 615 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 615, 'op': 'literal'}
    instructions[684] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 615 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 615, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[685] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 615 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 615, 'op': 'load'}
    instructions[686] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 615 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 615, 'op': 'add'}
    instructions[687] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 615 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 615, 'op': 'addl'}
    instructions[688] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 615 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 615, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[689] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 615 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 615, 'op': 'load'}
    instructions[690] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 615 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 615, 'op': 'store'}
    instructions[691] = {5'd0, 4'd8, 4'd0, 16'd18};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 616 {'literal': 18, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 616, 'op': 'literal'}
    instructions[692] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 616 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 616, 'op': 'store'}
    instructions[693] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 616 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 616, 'op': 'addl'}
    instructions[694] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 616 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 616, 'op': 'literal'}
    instructions[695] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 616 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 616, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[696] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 616 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 616, 'op': 'load'}
    instructions[697] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 616 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 616, 'op': 'add'}
    instructions[698] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 616 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 616, 'op': 'addl'}
    instructions[699] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 616 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 616, 'op': 'load'}
    instructions[700] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 616 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 616, 'op': 'store'}
    instructions[701] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 616 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 616, 'op': 'addl'}
    instructions[702] = {5'd0, 4'd8, 4'd0, 16'd608};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 616 {'literal': 608, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 616, 'op': 'literal'}
    instructions[703] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 616 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 616, 'op': 'store'}
    instructions[704] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 616 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 616, 'op': 'addl'}
    instructions[705] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 616 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 616, 'op': 'literal'}
    instructions[706] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 616 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 616, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[707] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 616 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 616, 'op': 'load'}
    instructions[708] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 616 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 616, 'op': 'add'}
    instructions[709] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 616 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 616, 'op': 'addl'}
    instructions[710] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 616 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 616, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[711] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 616 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 616, 'op': 'load'}
    instructions[712] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 616 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 616, 'op': 'store'}
    instructions[713] = {5'd0, 4'd8, 4'd0, 16'd18};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 617 {'literal': 18, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 617, 'op': 'literal'}
    instructions[714] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 617 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 617, 'op': 'store'}
    instructions[715] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 617 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 617, 'op': 'addl'}
    instructions[716] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 617 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 617, 'op': 'literal'}
    instructions[717] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 617 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 617, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[718] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 617 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 617, 'op': 'load'}
    instructions[719] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 617 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 617, 'op': 'add'}
    instructions[720] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 617 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 617, 'op': 'addl'}
    instructions[721] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 617 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 617, 'op': 'load'}
    instructions[722] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 617 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 617, 'op': 'store'}
    instructions[723] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 617 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 617, 'op': 'addl'}
    instructions[724] = {5'd0, 4'd8, 4'd0, 16'd14};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 617 {'literal': 14, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 617, 'op': 'literal'}
    instructions[725] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 617 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 617, 'op': 'store'}
    instructions[726] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 617 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 617, 'op': 'addl'}
    instructions[727] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 617 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 617, 'op': 'literal'}
    instructions[728] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 617 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 617, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[729] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 617 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 617, 'op': 'load'}
    instructions[730] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 617 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 617, 'op': 'add'}
    instructions[731] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 617 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 617, 'op': 'addl'}
    instructions[732] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 617 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 617, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[733] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 617 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 617, 'op': 'load'}
    instructions[734] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 617 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 617, 'op': 'store'}
    instructions[735] = {5'd0, 4'd8, 4'd0, 16'd18};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 618 {'literal': 18, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 618, 'op': 'literal'}
    instructions[736] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 618 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 618, 'op': 'store'}
    instructions[737] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 618 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 618, 'op': 'addl'}
    instructions[738] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 618 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 618, 'op': 'literal'}
    instructions[739] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 618 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 618, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[740] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 618 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 618, 'op': 'load'}
    instructions[741] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 618 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 618, 'op': 'add'}
    instructions[742] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 618 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 618, 'op': 'addl'}
    instructions[743] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 618 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 618, 'op': 'load'}
    instructions[744] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 618 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 618, 'op': 'store'}
    instructions[745] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 618 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 618, 'op': 'addl'}
    instructions[746] = {5'd0, 4'd8, 4'd0, 16'd14};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 618 {'literal': 14, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 618, 'op': 'literal'}
    instructions[747] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 618 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 618, 'op': 'store'}
    instructions[748] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 618 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 618, 'op': 'addl'}
    instructions[749] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 618 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 618, 'op': 'literal'}
    instructions[750] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 618 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 618, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[751] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 618 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 618, 'op': 'load'}
    instructions[752] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 618 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 618, 'op': 'add'}
    instructions[753] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 618 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 618, 'op': 'addl'}
    instructions[754] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 618 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 618, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[755] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 618 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 618, 'op': 'load'}
    instructions[756] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 618 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 618, 'op': 'store'}
    instructions[757] = {5'd0, 4'd8, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 619 {'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 619, 'op': 'literal'}
    instructions[758] = {5'd1, 4'd2, 4'd4, 16'd2062};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 619 {'a': 4, 'literal': 2062, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 619, 'op': 'addl'}
    instructions[759] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 619 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 619, 'op': 'store'}
    instructions[760] = {5'd10, 4'd0, 4'd0, 16'd761};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 614 {'label': 761, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 614, 'op': 'goto'}
    instructions[761] = {5'd10, 4'd0, 4'd0, 16'd907};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 621 {'label': 907, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 621, 'op': 'goto'}
    instructions[762] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625, 'op': 'store'}
    instructions[763] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625, 'op': 'addl'}
    instructions[764] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625, 'op': 'store'}
    instructions[765] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625, 'op': 'addl'}
    instructions[766] = {5'd0, 4'd8, 4'd0, 16'd561};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625 {'literal': 561, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625, 'op': 'literal'}
    instructions[767] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625, 'op': 'store'}
    instructions[768] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625, 'op': 'addl'}
    instructions[769] = {5'd0, 4'd8, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625 {'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625, 'op': 'literal'}
    instructions[770] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625, 'op': 'store'}
    instructions[771] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625, 'op': 'addl'}
    instructions[772] = {5'd0, 4'd8, 4'd0, 16'd581};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625 {'literal': 581, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625, 'op': 'literal'}
    instructions[773] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625, 'op': 'addl'}
    instructions[774] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625, 'op': 'load'}
    instructions[775] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625, 'op': 'store'}
    instructions[776] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625, 'op': 'addl'}
    instructions[777] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625, 'op': 'addl'}
    instructions[778] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625, 'op': 'addl'}
    instructions[779] = {5'd4, 4'd6, 4'd0, 16'd3325};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625 {'z': 6, 'label': 3325, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625, 'op': 'call'}
    instructions[780] = {5'd1, 4'd3, 4'd3, -16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625 {'a': 3, 'literal': -3, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625, 'op': 'addl'}
    instructions[781] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[782] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625, 'op': 'load'}
    instructions[783] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[784] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625, 'op': 'load'}
    instructions[785] = {5'd0, 4'd2, 4'd0, 16'd582};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625 {'literal': 582, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625, 'op': 'literal'}
    instructions[786] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625, 'op': 'load'}
    instructions[787] = {5'd1, 4'd2, 4'd4, 16'd2056};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625 {'a': 4, 'literal': 2056, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625, 'op': 'addl'}
    instructions[788] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 625, 'op': 'store'}
    instructions[789] = {5'd0, 4'd8, 4'd0, 16'd586};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 626 {'literal': 586, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 626, 'op': 'literal'}
    instructions[790] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 626 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 626, 'op': 'addl'}
    instructions[791] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 626 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 626, 'op': 'load'}
    instructions[792] = {5'd8, 4'd0, 4'd8, 16'd797};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 626 {'a': 8, 'label': 797, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 626, 'op': 'jmp_if_false'}
    instructions[793] = {5'd0, 4'd8, 4'd0, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 627 {'literal': 4, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 627, 'op': 'literal'}
    instructions[794] = {5'd1, 4'd2, 4'd4, 16'd2062};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 627 {'a': 4, 'literal': 2062, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 627, 'op': 'addl'}
    instructions[795] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 627 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 627, 'op': 'store'}
    instructions[796] = {5'd10, 4'd0, 4'd0, 16'd805};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 626 {'label': 805, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 626, 'op': 'goto'}
    instructions[797] = {5'd1, 4'd8, 4'd4, 16'd2051};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 628 {'a': 4, 'literal': 2051, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 628, 'op': 'addl'}
    instructions[798] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 628 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 628, 'op': 'addl'}
    instructions[799] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 628 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 628, 'op': 'load'}
    instructions[800] = {5'd8, 4'd0, 4'd8, 16'd805};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 628 {'a': 8, 'label': 805, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 628, 'op': 'jmp_if_false'}
    instructions[801] = {5'd0, 4'd8, 4'd0, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 629 {'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 629, 'op': 'literal'}
    instructions[802] = {5'd1, 4'd2, 4'd4, 16'd2062};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 629 {'a': 4, 'literal': 2062, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 629, 'op': 'addl'}
    instructions[803] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 629 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 629, 'op': 'store'}
    instructions[804] = {5'd10, 4'd0, 4'd0, 16'd805};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 628 {'label': 805, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 628, 'op': 'goto'}
    instructions[805] = {5'd10, 4'd0, 4'd0, 16'd907};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 631 {'label': 907, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 631, 'op': 'goto'}
    instructions[806] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636, 'op': 'store'}
    instructions[807] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636, 'op': 'addl'}
    instructions[808] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636, 'op': 'store'}
    instructions[809] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636, 'op': 'addl'}
    instructions[810] = {5'd0, 4'd8, 4'd0, 16'd561};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636 {'literal': 561, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636, 'op': 'literal'}
    instructions[811] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636, 'op': 'store'}
    instructions[812] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636, 'op': 'addl'}
    instructions[813] = {5'd0, 4'd8, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636 {'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636, 'op': 'literal'}
    instructions[814] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636, 'op': 'store'}
    instructions[815] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636, 'op': 'addl'}
    instructions[816] = {5'd0, 4'd8, 4'd0, 16'd581};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636 {'literal': 581, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636, 'op': 'literal'}
    instructions[817] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636, 'op': 'addl'}
    instructions[818] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636, 'op': 'load'}
    instructions[819] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636, 'op': 'store'}
    instructions[820] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636, 'op': 'addl'}
    instructions[821] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636, 'op': 'addl'}
    instructions[822] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636, 'op': 'addl'}
    instructions[823] = {5'd4, 4'd6, 4'd0, 16'd3325};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636 {'z': 6, 'label': 3325, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636, 'op': 'call'}
    instructions[824] = {5'd1, 4'd3, 4'd3, -16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636 {'a': 3, 'literal': -3, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636, 'op': 'addl'}
    instructions[825] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[826] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636, 'op': 'load'}
    instructions[827] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[828] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636, 'op': 'load'}
    instructions[829] = {5'd0, 4'd2, 4'd0, 16'd582};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636 {'literal': 582, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636, 'op': 'literal'}
    instructions[830] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636, 'op': 'load'}
    instructions[831] = {5'd1, 4'd2, 4'd4, 16'd2056};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636 {'a': 4, 'literal': 2056, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636, 'op': 'addl'}
    instructions[832] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 636, 'op': 'store'}
    instructions[833] = {5'd0, 4'd8, 4'd0, 16'd586};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 637 {'literal': 586, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 637, 'op': 'literal'}
    instructions[834] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 637 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 637, 'op': 'addl'}
    instructions[835] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 637 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 637, 'op': 'load'}
    instructions[836] = {5'd8, 4'd0, 4'd8, 16'd841};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 637 {'a': 8, 'label': 841, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 637, 'op': 'jmp_if_false'}
    instructions[837] = {5'd0, 4'd8, 4'd0, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 638 {'literal': 4, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 638, 'op': 'literal'}
    instructions[838] = {5'd1, 4'd2, 4'd4, 16'd2062};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 638 {'a': 4, 'literal': 2062, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 638, 'op': 'addl'}
    instructions[839] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 638 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 638, 'op': 'store'}
    instructions[840] = {5'd10, 4'd0, 4'd0, 16'd897};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 637 {'label': 897, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 637, 'op': 'goto'}
    instructions[841] = {5'd0, 4'd8, 4'd0, 16'd563};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 639 {'literal': 563, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 639, 'op': 'literal'}
    instructions[842] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 639 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 639, 'op': 'addl'}
    instructions[843] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 639 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 639, 'op': 'load'}
    instructions[844] = {5'd8, 4'd0, 4'd8, 16'd868};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640 {'a': 8, 'label': 868, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640, 'op': 'jmp_if_false'}
    instructions[845] = {5'd0, 4'd8, 4'd0, 16'd18};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640 {'literal': 18, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640, 'op': 'literal'}
    instructions[846] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640, 'op': 'store'}
    instructions[847] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640, 'op': 'addl'}
    instructions[848] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640, 'op': 'literal'}
    instructions[849] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[850] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640, 'op': 'load'}
    instructions[851] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640, 'op': 'add'}
    instructions[852] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640, 'op': 'addl'}
    instructions[853] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640, 'op': 'load'}
    instructions[854] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640, 'op': 'store'}
    instructions[855] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640, 'op': 'addl'}
    instructions[856] = {5'd0, 4'd8, 4'd0, 16'd14};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640 {'literal': 14, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640, 'op': 'literal'}
    instructions[857] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640, 'op': 'store'}
    instructions[858] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640, 'op': 'addl'}
    instructions[859] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640, 'op': 'literal'}
    instructions[860] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[861] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640, 'op': 'load'}
    instructions[862] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640, 'op': 'add'}
    instructions[863] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640, 'op': 'addl'}
    instructions[864] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640, 'op': 'load'}
    instructions[865] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[866] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640, 'op': 'load'}
    instructions[867] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 640, 'op': 'equal'}
    instructions[868] = {5'd8, 4'd0, 4'd8, 16'd892};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641 {'a': 8, 'label': 892, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641, 'op': 'jmp_if_false'}
    instructions[869] = {5'd0, 4'd8, 4'd0, 16'd18};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641 {'literal': 18, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641, 'op': 'literal'}
    instructions[870] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641, 'op': 'store'}
    instructions[871] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641, 'op': 'addl'}
    instructions[872] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641, 'op': 'literal'}
    instructions[873] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[874] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641, 'op': 'load'}
    instructions[875] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641, 'op': 'add'}
    instructions[876] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641, 'op': 'addl'}
    instructions[877] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641, 'op': 'load'}
    instructions[878] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641, 'op': 'store'}
    instructions[879] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641, 'op': 'addl'}
    instructions[880] = {5'd0, 4'd8, 4'd0, 16'd14};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641 {'literal': 14, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641, 'op': 'literal'}
    instructions[881] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641, 'op': 'store'}
    instructions[882] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641, 'op': 'addl'}
    instructions[883] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641, 'op': 'literal'}
    instructions[884] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[885] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641, 'op': 'load'}
    instructions[886] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641, 'op': 'add'}
    instructions[887] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641, 'op': 'addl'}
    instructions[888] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641, 'op': 'load'}
    instructions[889] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[890] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641, 'op': 'load'}
    instructions[891] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 641, 'op': 'equal'}
    instructions[892] = {5'd8, 4'd0, 4'd8, 16'd897};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 639 {'a': 8, 'label': 897, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 639, 'op': 'jmp_if_false'}
    instructions[893] = {5'd0, 4'd8, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 642 {'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 642, 'op': 'literal'}
    instructions[894] = {5'd1, 4'd2, 4'd4, 16'd2062};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 642 {'a': 4, 'literal': 2062, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 642, 'op': 'addl'}
    instructions[895] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 642 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 642, 'op': 'store'}
    instructions[896] = {5'd10, 4'd0, 4'd0, 16'd897};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 639 {'label': 897, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 639, 'op': 'goto'}
    instructions[897] = {5'd10, 4'd0, 4'd0, 16'd907};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 645 {'label': 907, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 645, 'op': 'goto'}
    instructions[898] = {5'd0, 4'd8, 4'd0, 16'd563};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 649 {'literal': 563, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 649, 'op': 'literal'}
    instructions[899] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 649 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 649, 'op': 'addl'}
    instructions[900] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 649 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 649, 'op': 'load'}
    instructions[901] = {5'd8, 4'd0, 4'd8, 16'd906};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 649 {'a': 8, 'label': 906, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 649, 'op': 'jmp_if_false'}
    instructions[902] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 649 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 649, 'op': 'literal'}
    instructions[903] = {5'd1, 4'd2, 4'd4, 16'd2062};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 649 {'a': 4, 'literal': 2062, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 649, 'op': 'addl'}
    instructions[904] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 649 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 649, 'op': 'store'}
    instructions[905] = {5'd10, 4'd0, 4'd0, 16'd906};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 649 {'label': 906, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 649, 'op': 'goto'}
    instructions[906] = {5'd10, 4'd0, 4'd0, 16'd907};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 650 {'label': 907, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 650, 'op': 'goto'}
    instructions[907] = {5'd0, 4'd8, 4'd0, 16'd587};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 653 {'literal': 587, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 653, 'op': 'literal'}
    instructions[908] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 653 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 653, 'op': 'addl'}
    instructions[909] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 653 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 653, 'op': 'load'}
    instructions[910] = {5'd8, 4'd0, 4'd8, 16'd915};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 653 {'a': 8, 'label': 915, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 653, 'op': 'jmp_if_false'}
    instructions[911] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 653 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 653, 'op': 'literal'}
    instructions[912] = {5'd1, 4'd2, 4'd4, 16'd2062};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 653 {'a': 4, 'literal': 2062, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 653, 'op': 'addl'}
    instructions[913] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 653 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 653, 'op': 'store'}
    instructions[914] = {5'd10, 4'd0, 4'd0, 16'd915};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 653 {'label': 915, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 653, 'op': 'goto'}
    instructions[915] = {5'd1, 4'd8, 4'd4, 16'd2056};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 656 {'a': 4, 'literal': 2056, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 656, 'op': 'addl'}
    instructions[916] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 656 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 656, 'op': 'addl'}
    instructions[917] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 656 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 656, 'op': 'load'}
    instructions[918] = {5'd8, 4'd0, 4'd8, 16'd980};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 656 {'a': 8, 'label': 980, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 656, 'op': 'jmp_if_false'}
    instructions[919] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657, 'op': 'store'}
    instructions[920] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657, 'op': 'addl'}
    instructions[921] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657, 'op': 'store'}
    instructions[922] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657, 'op': 'addl'}
    instructions[923] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657, 'op': 'addl'}
    instructions[924] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657, 'op': 'store'}
    instructions[925] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657, 'op': 'addl'}
    instructions[926] = {5'd0, 4'd8, 4'd0, 16'd21};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657 {'literal': 21, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657, 'op': 'literal'}
    instructions[927] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657, 'op': 'addl'}
    instructions[928] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657, 'op': 'load'}
    instructions[929] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657, 'op': 'store'}
    instructions[930] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657, 'op': 'addl'}
    instructions[931] = {5'd0, 4'd8, 4'd0, 16'd581};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657 {'literal': 581, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657, 'op': 'literal'}
    instructions[932] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657, 'op': 'addl'}
    instructions[933] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657, 'op': 'load'}
    instructions[934] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657, 'op': 'store'}
    instructions[935] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657, 'op': 'addl'}
    instructions[936] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657, 'op': 'addl'}
    instructions[937] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657, 'op': 'addl'}
    instructions[938] = {5'd4, 4'd6, 4'd0, 16'd5387};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657 {'z': 6, 'label': 5387, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657, 'op': 'call'}
    instructions[939] = {5'd1, 4'd3, 4'd3, -16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657 {'a': 3, 'literal': -3, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657, 'op': 'addl'}
    instructions[940] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[941] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657, 'op': 'load'}
    instructions[942] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[943] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657, 'op': 'load'}
    instructions[944] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 657, 'op': 'addl'}
    instructions[945] = {5'd1, 4'd8, 4'd4, 16'd2055};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659 {'a': 4, 'literal': 2055, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659, 'op': 'addl'}
    instructions[946] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659, 'op': 'addl'}
    instructions[947] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659, 'op': 'load'}
    instructions[948] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659, 'op': 'store'}
    instructions[949] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659, 'op': 'addl'}
    instructions[950] = {5'd1, 4'd8, 4'd4, 16'd2062};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659 {'a': 4, 'literal': 2062, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659, 'op': 'addl'}
    instructions[951] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659, 'op': 'addl'}
    instructions[952] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659, 'op': 'load'}
    instructions[953] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[954] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659, 'op': 'load'}
    instructions[955] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659, 'op': 'equal'}
    instructions[956] = {5'd8, 4'd0, 4'd8, 16'd979};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659 {'a': 8, 'label': 979, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659, 'op': 'jmp_if_false'}
    instructions[957] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659, 'op': 'store'}
    instructions[958] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659, 'op': 'addl'}
    instructions[959] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659, 'op': 'store'}
    instructions[960] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659, 'op': 'addl'}
    instructions[961] = {5'd1, 4'd8, 4'd4, 16'd1024};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659 {'a': 4, 'literal': 1024, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659, 'op': 'addl'}
    instructions[962] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659, 'op': 'store'}
    instructions[963] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659, 'op': 'addl'}
    instructions[964] = {5'd1, 4'd8, 4'd4, 16'd2051};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659 {'a': 4, 'literal': 2051, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659, 'op': 'addl'}
    instructions[965] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659, 'op': 'addl'}
    instructions[966] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659, 'op': 'load'}
    instructions[967] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659, 'op': 'store'}
    instructions[968] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659, 'op': 'addl'}
    instructions[969] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659, 'op': 'addl'}
    instructions[970] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659, 'op': 'addl'}
    instructions[971] = {5'd4, 4'd6, 4'd0, 16'd1040};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659 {'z': 6, 'label': 1040, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659, 'op': 'call'}
    instructions[972] = {5'd1, 4'd3, 4'd3, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659 {'a': 3, 'literal': -2, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659, 'op': 'addl'}
    instructions[973] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[974] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659, 'op': 'load'}
    instructions[975] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[976] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659, 'op': 'load'}
    instructions[977] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659, 'op': 'addl'}
    instructions[978] = {5'd10, 4'd0, 4'd0, 16'd979};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659 {'label': 979, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 659, 'op': 'goto'}
    instructions[979] = {5'd10, 4'd0, 4'd0, 16'd980};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 656 {'label': 980, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 656, 'op': 'goto'}
    instructions[980] = {5'd0, 4'd8, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 662 {'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 662, 'op': 'literal'}
    instructions[981] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 662 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 662, 'op': 'store'}
    instructions[982] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 662 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 662, 'op': 'addl'}
    instructions[983] = {5'd1, 4'd8, 4'd4, 16'd2062};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 662 {'a': 4, 'literal': 2062, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 662, 'op': 'addl'}
    instructions[984] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 662 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 662, 'op': 'addl'}
    instructions[985] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 662 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 662, 'op': 'load'}
    instructions[986] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 662 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 662, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[987] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 662 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 662, 'op': 'load'}
    instructions[988] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 662 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 662, 'op': 'equal'}
    instructions[989] = {5'd8, 4'd0, 4'd8, 16'd994};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 662 {'a': 8, 'label': 994, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 662, 'op': 'jmp_if_false'}
    instructions[990] = {5'd0, 4'd8, 4'd0, 16'd16};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 662 {'literal': 16, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 662, 'op': 'literal'}
    instructions[991] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 662 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 662, 'op': 'addl'}
    instructions[992] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 662 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 662, 'op': 'load'}
    instructions[993] = {5'd14, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 662 {'a': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 662, 'op': 'ready'}
    instructions[994] = {5'd8, 4'd0, 4'd8, 16'd997};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 662 {'a': 8, 'label': 997, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 662, 'op': 'jmp_if_false'}
    instructions[995] = {5'd10, 4'd0, 4'd0, 16'd1036};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 663 {'label': 1036, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 663, 'op': 'goto'}
    instructions[996] = {5'd10, 4'd0, 4'd0, 16'd997};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 662 {'label': 997, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 662, 'op': 'goto'}
    instructions[997] = {5'd1, 4'd8, 4'd4, 16'd2055};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 666 {'a': 4, 'literal': 2055, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 666, 'op': 'addl'}
    instructions[998] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 666 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 666, 'op': 'addl'}
    instructions[999] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 666 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 666, 'op': 'load'}
    instructions[1000] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 666 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 666, 'op': 'store'}
    instructions[1001] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 666 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 666, 'op': 'addl'}
    instructions[1002] = {5'd1, 4'd8, 4'd4, 16'd2062};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 666 {'a': 4, 'literal': 2062, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 666, 'op': 'addl'}
    instructions[1003] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 666 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 666, 'op': 'addl'}
    instructions[1004] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 666 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 666, 'op': 'load'}
    instructions[1005] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 666 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 666, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1006] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 666 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 666, 'op': 'load'}
    instructions[1007] = {5'd13, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 666 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 666, 'op': 'not_equal'}
    instructions[1008] = {5'd8, 4'd0, 4'd8, 16'd1014};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 666 {'a': 8, 'label': 1014, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 666, 'op': 'jmp_if_false'}
    instructions[1009] = {5'd0, 4'd8, 4'd0, 16'd120};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 667 {'literal': 120, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 667, 'op': 'literal'}
    instructions[1010] = {5'd1, 4'd2, 4'd4, 16'd2052};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 667 {'a': 4, 'literal': 2052, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 667, 'op': 'addl'}
    instructions[1011] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 667 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 667, 'op': 'store'}
    instructions[1012] = {5'd10, 4'd0, 4'd0, 16'd1036};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 668 {'label': 1036, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 668, 'op': 'goto'}
    instructions[1013] = {5'd10, 4'd0, 4'd0, 16'd1014};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 666 {'label': 1014, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 666, 'op': 'goto'}
    instructions[1014] = {5'd10, 4'd0, 4'd0, 16'd1017};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 596 {'label': 1017, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 596, 'op': 'goto'}
    instructions[1015] = {5'd0, 4'd8, 4'd0, 16'd1000};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 672 {'literal': 1000, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 672, 'op': 'literal'}
    instructions[1016] = {5'd15, 4'd0, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 672 {'a': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 672, 'op': 'wait_clocks'}
    instructions[1017] = {5'd1, 4'd8, 4'd4, 16'd2053};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594 {'a': 4, 'literal': 2053, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594, 'op': 'addl'}
    instructions[1018] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594, 'op': 'addl'}
    instructions[1019] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594, 'op': 'load'}
    instructions[1020] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594, 'op': 'store'}
    instructions[1021] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594, 'op': 'addl'}
    instructions[1022] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594, 'op': 'literal'}
    instructions[1023] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594, 'op': 'store'}
    instructions[1024] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594, 'op': 'addl'}
    instructions[1025] = {5'd1, 4'd8, 4'd4, 16'd2053};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594 {'a': 4, 'literal': 2053, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594, 'op': 'addl'}
    instructions[1026] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594, 'op': 'addl'}
    instructions[1027] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594, 'op': 'load'}
    instructions[1028] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1029] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594, 'op': 'load'}
    instructions[1030] = {5'd9, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594, 'op': 'subtract'}
    instructions[1031] = {5'd1, 4'd2, 4'd4, 16'd2053};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594 {'a': 4, 'literal': 2053, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594, 'op': 'addl'}
    instructions[1032] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594, 'op': 'store'}
    instructions[1033] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1034] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594, 'op': 'load'}
    instructions[1035] = {5'd10, 4'd0, 4'd0, 16'd546};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594 {'label': 546, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 594, 'op': 'goto'}
    instructions[1036] = {5'd10, 4'd0, 4'd0, 16'd180};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 536 {'label': 180, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 536, 'op': 'goto'}
    instructions[1037] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 508 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 508, 'op': 'addl'}
    instructions[1038] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 508 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 508, 'op': 'addl'}
    instructions[1039] = {5'd16, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 508 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 508, 'op': 'return'}
    instructions[1040] = {5'd1, 4'd3, 4'd3, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 389 {'a': 3, 'literal': 4, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 389, 'op': 'addl'}
    instructions[1041] = {5'd0, 4'd8, 4'd0, 16'd17};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 391 {'literal': 17, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 391, 'op': 'literal'}
    instructions[1042] = {5'd1, 4'd2, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 391 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 391, 'op': 'addl'}
    instructions[1043] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 391 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 391, 'op': 'store'}
    instructions[1044] = {5'd0, 4'd8, 4'd0, 16'd610};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397 {'literal': 610, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397, 'op': 'literal'}
    instructions[1045] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397, 'op': 'addl'}
    instructions[1046] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397, 'op': 'load'}
    instructions[1047] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397, 'op': 'store'}
    instructions[1048] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397, 'op': 'addl'}
    instructions[1049] = {5'd1, 4'd8, 4'd4, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397 {'a': 4, 'literal': -2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397, 'op': 'addl'}
    instructions[1050] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397, 'op': 'addl'}
    instructions[1051] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397, 'op': 'load'}
    instructions[1052] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397, 'op': 'store'}
    instructions[1053] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397, 'op': 'addl'}
    instructions[1054] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397, 'op': 'literal'}
    instructions[1055] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397, 'op': 'store'}
    instructions[1056] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397, 'op': 'addl'}
    instructions[1057] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397, 'op': 'addl'}
    instructions[1058] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397, 'op': 'addl'}
    instructions[1059] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397, 'op': 'load'}
    instructions[1060] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1061] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397, 'op': 'load'}
    instructions[1062] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397, 'op': 'add'}
    instructions[1063] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1064] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397, 'op': 'load'}
    instructions[1065] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397, 'op': 'add'}
    instructions[1066] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397, 'op': 'addl'}
    instructions[1067] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1068] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397, 'op': 'load'}
    instructions[1069] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 397, 'op': 'store'}
    instructions[1070] = {5'd0, 4'd8, 4'd0, 16'd23};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398 {'literal': 23, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398, 'op': 'literal'}
    instructions[1071] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398, 'op': 'addl'}
    instructions[1072] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398, 'op': 'load'}
    instructions[1073] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398, 'op': 'store'}
    instructions[1074] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398, 'op': 'addl'}
    instructions[1075] = {5'd1, 4'd8, 4'd4, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398 {'a': 4, 'literal': -2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398, 'op': 'addl'}
    instructions[1076] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398, 'op': 'addl'}
    instructions[1077] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398, 'op': 'load'}
    instructions[1078] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398, 'op': 'store'}
    instructions[1079] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398, 'op': 'addl'}
    instructions[1080] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398, 'op': 'literal'}
    instructions[1081] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398, 'op': 'store'}
    instructions[1082] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398, 'op': 'addl'}
    instructions[1083] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398, 'op': 'addl'}
    instructions[1084] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398, 'op': 'addl'}
    instructions[1085] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398, 'op': 'load'}
    instructions[1086] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1087] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398, 'op': 'load'}
    instructions[1088] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398, 'op': 'add'}
    instructions[1089] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1090] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398, 'op': 'load'}
    instructions[1091] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398, 'op': 'add'}
    instructions[1092] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398, 'op': 'addl'}
    instructions[1093] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1094] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398, 'op': 'load'}
    instructions[1095] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 398, 'op': 'store'}
    instructions[1096] = {5'd0, 4'd8, 4'd0, 16'd608};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399 {'literal': 608, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399, 'op': 'literal'}
    instructions[1097] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399, 'op': 'store'}
    instructions[1098] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399, 'op': 'addl'}
    instructions[1099] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399, 'op': 'literal'}
    instructions[1100] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1101] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399, 'op': 'load'}
    instructions[1102] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399, 'op': 'add'}
    instructions[1103] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399, 'op': 'addl'}
    instructions[1104] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399, 'op': 'load'}
    instructions[1105] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399, 'op': 'store'}
    instructions[1106] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399, 'op': 'addl'}
    instructions[1107] = {5'd1, 4'd8, 4'd4, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399 {'a': 4, 'literal': -2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399, 'op': 'addl'}
    instructions[1108] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399, 'op': 'addl'}
    instructions[1109] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399, 'op': 'load'}
    instructions[1110] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399, 'op': 'store'}
    instructions[1111] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399, 'op': 'addl'}
    instructions[1112] = {5'd0, 4'd8, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399 {'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399, 'op': 'literal'}
    instructions[1113] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399, 'op': 'store'}
    instructions[1114] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399, 'op': 'addl'}
    instructions[1115] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399, 'op': 'addl'}
    instructions[1116] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399, 'op': 'addl'}
    instructions[1117] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399, 'op': 'load'}
    instructions[1118] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1119] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399, 'op': 'load'}
    instructions[1120] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399, 'op': 'add'}
    instructions[1121] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1122] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399, 'op': 'load'}
    instructions[1123] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399, 'op': 'add'}
    instructions[1124] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399, 'op': 'addl'}
    instructions[1125] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1126] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399, 'op': 'load'}
    instructions[1127] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 399, 'op': 'store'}
    instructions[1128] = {5'd0, 4'd8, 4'd0, 16'd608};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400 {'literal': 608, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400, 'op': 'literal'}
    instructions[1129] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400, 'op': 'store'}
    instructions[1130] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400, 'op': 'addl'}
    instructions[1131] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400, 'op': 'literal'}
    instructions[1132] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1133] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400, 'op': 'load'}
    instructions[1134] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400, 'op': 'add'}
    instructions[1135] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400, 'op': 'addl'}
    instructions[1136] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400, 'op': 'load'}
    instructions[1137] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400, 'op': 'store'}
    instructions[1138] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400, 'op': 'addl'}
    instructions[1139] = {5'd1, 4'd8, 4'd4, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400 {'a': 4, 'literal': -2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400, 'op': 'addl'}
    instructions[1140] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400, 'op': 'addl'}
    instructions[1141] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400, 'op': 'load'}
    instructions[1142] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400, 'op': 'store'}
    instructions[1143] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400, 'op': 'addl'}
    instructions[1144] = {5'd0, 4'd8, 4'd0, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400 {'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400, 'op': 'literal'}
    instructions[1145] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400, 'op': 'store'}
    instructions[1146] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400, 'op': 'addl'}
    instructions[1147] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400, 'op': 'addl'}
    instructions[1148] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400, 'op': 'addl'}
    instructions[1149] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400, 'op': 'load'}
    instructions[1150] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1151] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400, 'op': 'load'}
    instructions[1152] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400, 'op': 'add'}
    instructions[1153] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1154] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400, 'op': 'load'}
    instructions[1155] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400, 'op': 'add'}
    instructions[1156] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400, 'op': 'addl'}
    instructions[1157] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1158] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400, 'op': 'load'}
    instructions[1159] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 400, 'op': 'store'}
    instructions[1160] = {5'd0, 4'd8, 4'd0, 16'd561};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401 {'literal': 561, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401, 'op': 'literal'}
    instructions[1161] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401, 'op': 'store'}
    instructions[1162] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401, 'op': 'addl'}
    instructions[1163] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401, 'op': 'literal'}
    instructions[1164] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1165] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401, 'op': 'load'}
    instructions[1166] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401, 'op': 'add'}
    instructions[1167] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401, 'op': 'addl'}
    instructions[1168] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401, 'op': 'load'}
    instructions[1169] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401, 'op': 'store'}
    instructions[1170] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401, 'op': 'addl'}
    instructions[1171] = {5'd1, 4'd8, 4'd4, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401 {'a': 4, 'literal': -2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401, 'op': 'addl'}
    instructions[1172] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401, 'op': 'addl'}
    instructions[1173] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401, 'op': 'load'}
    instructions[1174] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401, 'op': 'store'}
    instructions[1175] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401, 'op': 'addl'}
    instructions[1176] = {5'd0, 4'd8, 4'd0, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401 {'literal': 4, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401, 'op': 'literal'}
    instructions[1177] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401, 'op': 'store'}
    instructions[1178] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401, 'op': 'addl'}
    instructions[1179] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401, 'op': 'addl'}
    instructions[1180] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401, 'op': 'addl'}
    instructions[1181] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401, 'op': 'load'}
    instructions[1182] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1183] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401, 'op': 'load'}
    instructions[1184] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401, 'op': 'add'}
    instructions[1185] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1186] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401, 'op': 'load'}
    instructions[1187] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401, 'op': 'add'}
    instructions[1188] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401, 'op': 'addl'}
    instructions[1189] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1190] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401, 'op': 'load'}
    instructions[1191] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 401, 'op': 'store'}
    instructions[1192] = {5'd0, 4'd8, 4'd0, 16'd561};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402 {'literal': 561, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402, 'op': 'literal'}
    instructions[1193] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402, 'op': 'store'}
    instructions[1194] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402, 'op': 'addl'}
    instructions[1195] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402, 'op': 'literal'}
    instructions[1196] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1197] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402, 'op': 'load'}
    instructions[1198] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402, 'op': 'add'}
    instructions[1199] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402, 'op': 'addl'}
    instructions[1200] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402, 'op': 'load'}
    instructions[1201] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402, 'op': 'store'}
    instructions[1202] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402, 'op': 'addl'}
    instructions[1203] = {5'd1, 4'd8, 4'd4, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402 {'a': 4, 'literal': -2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402, 'op': 'addl'}
    instructions[1204] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402, 'op': 'addl'}
    instructions[1205] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402, 'op': 'load'}
    instructions[1206] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402, 'op': 'store'}
    instructions[1207] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402, 'op': 'addl'}
    instructions[1208] = {5'd0, 4'd8, 4'd0, 16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402 {'literal': 5, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402, 'op': 'literal'}
    instructions[1209] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402, 'op': 'store'}
    instructions[1210] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402, 'op': 'addl'}
    instructions[1211] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402, 'op': 'addl'}
    instructions[1212] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402, 'op': 'addl'}
    instructions[1213] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402, 'op': 'load'}
    instructions[1214] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1215] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402, 'op': 'load'}
    instructions[1216] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402, 'op': 'add'}
    instructions[1217] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1218] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402, 'op': 'load'}
    instructions[1219] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402, 'op': 'add'}
    instructions[1220] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402, 'op': 'addl'}
    instructions[1221] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1222] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402, 'op': 'load'}
    instructions[1223] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 402, 'op': 'store'}
    instructions[1224] = {5'd0, 4'd8, 4'd0, 16'd20480};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403 {'literal': 20480, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403, 'op': 'literal'}
    instructions[1225] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403, 'op': 'store'}
    instructions[1226] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403, 'op': 'addl'}
    instructions[1227] = {5'd1, 4'd8, 4'd4, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403 {'a': 4, 'literal': -2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403, 'op': 'addl'}
    instructions[1228] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403, 'op': 'addl'}
    instructions[1229] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403, 'op': 'load'}
    instructions[1230] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403, 'op': 'store'}
    instructions[1231] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403, 'op': 'addl'}
    instructions[1232] = {5'd0, 4'd8, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403 {'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403, 'op': 'literal'}
    instructions[1233] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403, 'op': 'store'}
    instructions[1234] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403, 'op': 'addl'}
    instructions[1235] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403, 'op': 'addl'}
    instructions[1236] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403, 'op': 'addl'}
    instructions[1237] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403, 'op': 'load'}
    instructions[1238] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1239] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403, 'op': 'load'}
    instructions[1240] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403, 'op': 'add'}
    instructions[1241] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1242] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403, 'op': 'load'}
    instructions[1243] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403, 'op': 'add'}
    instructions[1244] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403, 'op': 'addl'}
    instructions[1245] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1246] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403, 'op': 'load'}
    instructions[1247] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 403, 'op': 'store'}
    instructions[1248] = {5'd0, 4'd8, 4'd0, 16'd653};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404 {'literal': 653, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404, 'op': 'literal'}
    instructions[1249] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404, 'op': 'addl'}
    instructions[1250] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404, 'op': 'load'}
    instructions[1251] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404, 'op': 'store'}
    instructions[1252] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404, 'op': 'addl'}
    instructions[1253] = {5'd1, 4'd8, 4'd4, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404 {'a': 4, 'literal': -2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404, 'op': 'addl'}
    instructions[1254] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404, 'op': 'addl'}
    instructions[1255] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404, 'op': 'load'}
    instructions[1256] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404, 'op': 'store'}
    instructions[1257] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404, 'op': 'addl'}
    instructions[1258] = {5'd0, 4'd8, 4'd0, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404 {'literal': 7, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404, 'op': 'literal'}
    instructions[1259] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404, 'op': 'store'}
    instructions[1260] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404, 'op': 'addl'}
    instructions[1261] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404, 'op': 'addl'}
    instructions[1262] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404, 'op': 'addl'}
    instructions[1263] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404, 'op': 'load'}
    instructions[1264] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1265] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404, 'op': 'load'}
    instructions[1266] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404, 'op': 'add'}
    instructions[1267] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1268] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404, 'op': 'load'}
    instructions[1269] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404, 'op': 'add'}
    instructions[1270] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404, 'op': 'addl'}
    instructions[1271] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1272] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404, 'op': 'load'}
    instructions[1273] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 404, 'op': 'store'}
    instructions[1274] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405, 'op': 'literal'}
    instructions[1275] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405, 'op': 'store'}
    instructions[1276] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405, 'op': 'addl'}
    instructions[1277] = {5'd1, 4'd8, 4'd4, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405 {'a': 4, 'literal': -2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405, 'op': 'addl'}
    instructions[1278] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405, 'op': 'addl'}
    instructions[1279] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405, 'op': 'load'}
    instructions[1280] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405, 'op': 'store'}
    instructions[1281] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405, 'op': 'addl'}
    instructions[1282] = {5'd0, 4'd8, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405 {'literal': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405, 'op': 'literal'}
    instructions[1283] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405, 'op': 'store'}
    instructions[1284] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405, 'op': 'addl'}
    instructions[1285] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405, 'op': 'addl'}
    instructions[1286] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405, 'op': 'addl'}
    instructions[1287] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405, 'op': 'load'}
    instructions[1288] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1289] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405, 'op': 'load'}
    instructions[1290] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405, 'op': 'add'}
    instructions[1291] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1292] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405, 'op': 'load'}
    instructions[1293] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405, 'op': 'add'}
    instructions[1294] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405, 'op': 'addl'}
    instructions[1295] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1296] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405, 'op': 'load'}
    instructions[1297] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 405, 'op': 'store'}
    instructions[1298] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406, 'op': 'literal'}
    instructions[1299] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406, 'op': 'store'}
    instructions[1300] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406, 'op': 'addl'}
    instructions[1301] = {5'd1, 4'd8, 4'd4, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406 {'a': 4, 'literal': -2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406, 'op': 'addl'}
    instructions[1302] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406, 'op': 'addl'}
    instructions[1303] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406, 'op': 'load'}
    instructions[1304] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406, 'op': 'store'}
    instructions[1305] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406, 'op': 'addl'}
    instructions[1306] = {5'd0, 4'd8, 4'd0, 16'd9};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406 {'literal': 9, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406, 'op': 'literal'}
    instructions[1307] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406, 'op': 'store'}
    instructions[1308] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406, 'op': 'addl'}
    instructions[1309] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406, 'op': 'addl'}
    instructions[1310] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406, 'op': 'addl'}
    instructions[1311] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406, 'op': 'load'}
    instructions[1312] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1313] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406, 'op': 'load'}
    instructions[1314] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406, 'op': 'add'}
    instructions[1315] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1316] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406, 'op': 'load'}
    instructions[1317] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406, 'op': 'add'}
    instructions[1318] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406, 'op': 'addl'}
    instructions[1319] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1320] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406, 'op': 'load'}
    instructions[1321] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 406, 'op': 'store'}
    instructions[1322] = {5'd0, 4'd8, 4'd0, 16'd12};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'literal': 12, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'op': 'literal'}
    instructions[1323] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'op': 'addl'}
    instructions[1324] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'op': 'load'}
    instructions[1325] = {5'd8, 4'd0, 4'd8, 16'd1375};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 8, 'label': 1375, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'op': 'jmp_if_false'}
    instructions[1326] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'op': 'literal'}
    instructions[1327] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'op': 'store'}
    instructions[1328] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'op': 'addl'}
    instructions[1329] = {5'd1, 4'd8, 4'd4, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 4, 'literal': -2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'op': 'addl'}
    instructions[1330] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'op': 'addl'}
    instructions[1331] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'op': 'load'}
    instructions[1332] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'op': 'store'}
    instructions[1333] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'op': 'addl'}
    instructions[1334] = {5'd0, 4'd8, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'op': 'literal'}
    instructions[1335] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'op': 'store'}
    instructions[1336] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'op': 'addl'}
    instructions[1337] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'op': 'addl'}
    instructions[1338] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'op': 'addl'}
    instructions[1339] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'op': 'load'}
    instructions[1340] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1341] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'op': 'load'}
    instructions[1342] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'op': 'add'}
    instructions[1343] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1344] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'op': 'load'}
    instructions[1345] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'op': 'add'}
    instructions[1346] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'op': 'addl'}
    instructions[1347] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'op': 'load'}
    instructions[1348] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1349] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'op': 'load'}
    instructions[1350] = {5'd17, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'op': 'or'}
    instructions[1351] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'op': 'store'}
    instructions[1352] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'op': 'addl'}
    instructions[1353] = {5'd1, 4'd8, 4'd4, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 4, 'literal': -2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'op': 'addl'}
    instructions[1354] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'op': 'addl'}
    instructions[1355] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'op': 'load'}
    instructions[1356] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'op': 'store'}
    instructions[1357] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'op': 'addl'}
    instructions[1358] = {5'd0, 4'd8, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'op': 'literal'}
    instructions[1359] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'op': 'store'}
    instructions[1360] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'op': 'addl'}
    instructions[1361] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'op': 'addl'}
    instructions[1362] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'op': 'addl'}
    instructions[1363] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'op': 'load'}
    instructions[1364] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1365] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'op': 'load'}
    instructions[1366] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'op': 'add'}
    instructions[1367] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1368] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'op': 'load'}
    instructions[1369] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'op': 'add'}
    instructions[1370] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'op': 'addl'}
    instructions[1371] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1372] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'op': 'load'}
    instructions[1373] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'op': 'store'}
    instructions[1374] = {5'd10, 4'd0, 4'd0, 16'd1375};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409 {'label': 1375, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 409, 'op': 'goto'}
    instructions[1375] = {5'd0, 4'd8, 4'd0, 16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'literal': 5, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'op': 'literal'}
    instructions[1376] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'op': 'addl'}
    instructions[1377] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'op': 'load'}
    instructions[1378] = {5'd8, 4'd0, 4'd8, 16'd1428};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 8, 'label': 1428, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'op': 'jmp_if_false'}
    instructions[1379] = {5'd0, 4'd8, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'op': 'literal'}
    instructions[1380] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'op': 'store'}
    instructions[1381] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'op': 'addl'}
    instructions[1382] = {5'd1, 4'd8, 4'd4, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 4, 'literal': -2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'op': 'addl'}
    instructions[1383] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'op': 'addl'}
    instructions[1384] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'op': 'load'}
    instructions[1385] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'op': 'store'}
    instructions[1386] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'op': 'addl'}
    instructions[1387] = {5'd0, 4'd8, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'op': 'literal'}
    instructions[1388] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'op': 'store'}
    instructions[1389] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'op': 'addl'}
    instructions[1390] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'op': 'addl'}
    instructions[1391] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'op': 'addl'}
    instructions[1392] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'op': 'load'}
    instructions[1393] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1394] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'op': 'load'}
    instructions[1395] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'op': 'add'}
    instructions[1396] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1397] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'op': 'load'}
    instructions[1398] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'op': 'add'}
    instructions[1399] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'op': 'addl'}
    instructions[1400] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'op': 'load'}
    instructions[1401] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1402] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'op': 'load'}
    instructions[1403] = {5'd17, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'op': 'or'}
    instructions[1404] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'op': 'store'}
    instructions[1405] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'op': 'addl'}
    instructions[1406] = {5'd1, 4'd8, 4'd4, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 4, 'literal': -2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'op': 'addl'}
    instructions[1407] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'op': 'addl'}
    instructions[1408] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'op': 'load'}
    instructions[1409] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'op': 'store'}
    instructions[1410] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'op': 'addl'}
    instructions[1411] = {5'd0, 4'd8, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'op': 'literal'}
    instructions[1412] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'op': 'store'}
    instructions[1413] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'op': 'addl'}
    instructions[1414] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'op': 'addl'}
    instructions[1415] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'op': 'addl'}
    instructions[1416] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'op': 'load'}
    instructions[1417] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1418] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'op': 'load'}
    instructions[1419] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'op': 'add'}
    instructions[1420] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1421] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'op': 'load'}
    instructions[1422] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'op': 'add'}
    instructions[1423] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'op': 'addl'}
    instructions[1424] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1425] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'op': 'load'}
    instructions[1426] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'op': 'store'}
    instructions[1427] = {5'd10, 4'd0, 4'd0, 16'd1428};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410 {'label': 1428, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 410, 'op': 'goto'}
    instructions[1428] = {5'd0, 4'd8, 4'd0, 16'd22};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'literal': 22, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'op': 'literal'}
    instructions[1429] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'op': 'addl'}
    instructions[1430] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'op': 'load'}
    instructions[1431] = {5'd8, 4'd0, 4'd8, 16'd1481};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 8, 'label': 1481, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'op': 'jmp_if_false'}
    instructions[1432] = {5'd0, 4'd8, 4'd0, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'literal': 4, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'op': 'literal'}
    instructions[1433] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'op': 'store'}
    instructions[1434] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'op': 'addl'}
    instructions[1435] = {5'd1, 4'd8, 4'd4, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 4, 'literal': -2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'op': 'addl'}
    instructions[1436] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'op': 'addl'}
    instructions[1437] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'op': 'load'}
    instructions[1438] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'op': 'store'}
    instructions[1439] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'op': 'addl'}
    instructions[1440] = {5'd0, 4'd8, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'op': 'literal'}
    instructions[1441] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'op': 'store'}
    instructions[1442] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'op': 'addl'}
    instructions[1443] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'op': 'addl'}
    instructions[1444] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'op': 'addl'}
    instructions[1445] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'op': 'load'}
    instructions[1446] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1447] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'op': 'load'}
    instructions[1448] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'op': 'add'}
    instructions[1449] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1450] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'op': 'load'}
    instructions[1451] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'op': 'add'}
    instructions[1452] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'op': 'addl'}
    instructions[1453] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'op': 'load'}
    instructions[1454] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1455] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'op': 'load'}
    instructions[1456] = {5'd17, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'op': 'or'}
    instructions[1457] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'op': 'store'}
    instructions[1458] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'op': 'addl'}
    instructions[1459] = {5'd1, 4'd8, 4'd4, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 4, 'literal': -2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'op': 'addl'}
    instructions[1460] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'op': 'addl'}
    instructions[1461] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'op': 'load'}
    instructions[1462] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'op': 'store'}
    instructions[1463] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'op': 'addl'}
    instructions[1464] = {5'd0, 4'd8, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'op': 'literal'}
    instructions[1465] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'op': 'store'}
    instructions[1466] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'op': 'addl'}
    instructions[1467] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'op': 'addl'}
    instructions[1468] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'op': 'addl'}
    instructions[1469] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'op': 'load'}
    instructions[1470] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1471] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'op': 'load'}
    instructions[1472] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'op': 'add'}
    instructions[1473] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1474] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'op': 'load'}
    instructions[1475] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'op': 'add'}
    instructions[1476] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'op': 'addl'}
    instructions[1477] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1478] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'op': 'load'}
    instructions[1479] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'op': 'store'}
    instructions[1480] = {5'd10, 4'd0, 4'd0, 16'd1481};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411 {'label': 1481, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 411, 'op': 'goto'}
    instructions[1481] = {5'd0, 4'd8, 4'd0, 16'd649};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'literal': 649, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'op': 'literal'}
    instructions[1482] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'op': 'addl'}
    instructions[1483] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'op': 'load'}
    instructions[1484] = {5'd8, 4'd0, 4'd8, 16'd1534};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 8, 'label': 1534, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'op': 'jmp_if_false'}
    instructions[1485] = {5'd0, 4'd8, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'literal': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'op': 'literal'}
    instructions[1486] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'op': 'store'}
    instructions[1487] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'op': 'addl'}
    instructions[1488] = {5'd1, 4'd8, 4'd4, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 4, 'literal': -2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'op': 'addl'}
    instructions[1489] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'op': 'addl'}
    instructions[1490] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'op': 'load'}
    instructions[1491] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'op': 'store'}
    instructions[1492] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'op': 'addl'}
    instructions[1493] = {5'd0, 4'd8, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'op': 'literal'}
    instructions[1494] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'op': 'store'}
    instructions[1495] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'op': 'addl'}
    instructions[1496] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'op': 'addl'}
    instructions[1497] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'op': 'addl'}
    instructions[1498] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'op': 'load'}
    instructions[1499] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1500] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'op': 'load'}
    instructions[1501] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'op': 'add'}
    instructions[1502] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1503] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'op': 'load'}
    instructions[1504] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'op': 'add'}
    instructions[1505] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'op': 'addl'}
    instructions[1506] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'op': 'load'}
    instructions[1507] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1508] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'op': 'load'}
    instructions[1509] = {5'd17, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'op': 'or'}
    instructions[1510] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'op': 'store'}
    instructions[1511] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'op': 'addl'}
    instructions[1512] = {5'd1, 4'd8, 4'd4, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 4, 'literal': -2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'op': 'addl'}
    instructions[1513] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'op': 'addl'}
    instructions[1514] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'op': 'load'}
    instructions[1515] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'op': 'store'}
    instructions[1516] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'op': 'addl'}
    instructions[1517] = {5'd0, 4'd8, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'op': 'literal'}
    instructions[1518] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'op': 'store'}
    instructions[1519] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'op': 'addl'}
    instructions[1520] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'op': 'addl'}
    instructions[1521] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'op': 'addl'}
    instructions[1522] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'op': 'load'}
    instructions[1523] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1524] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'op': 'load'}
    instructions[1525] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'op': 'add'}
    instructions[1526] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1527] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'op': 'load'}
    instructions[1528] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'op': 'add'}
    instructions[1529] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'op': 'addl'}
    instructions[1530] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1531] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'op': 'load'}
    instructions[1532] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'op': 'store'}
    instructions[1533] = {5'd10, 4'd0, 4'd0, 16'd1534};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412 {'label': 1534, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 412, 'op': 'goto'}
    instructions[1534] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'op': 'literal'}
    instructions[1535] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'op': 'addl'}
    instructions[1536] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'op': 'load'}
    instructions[1537] = {5'd8, 4'd0, 4'd8, 16'd1587};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 8, 'label': 1587, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'op': 'jmp_if_false'}
    instructions[1538] = {5'd0, 4'd8, 4'd0, 16'd16};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'literal': 16, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'op': 'literal'}
    instructions[1539] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'op': 'store'}
    instructions[1540] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'op': 'addl'}
    instructions[1541] = {5'd1, 4'd8, 4'd4, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 4, 'literal': -2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'op': 'addl'}
    instructions[1542] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'op': 'addl'}
    instructions[1543] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'op': 'load'}
    instructions[1544] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'op': 'store'}
    instructions[1545] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'op': 'addl'}
    instructions[1546] = {5'd0, 4'd8, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'op': 'literal'}
    instructions[1547] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'op': 'store'}
    instructions[1548] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'op': 'addl'}
    instructions[1549] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'op': 'addl'}
    instructions[1550] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'op': 'addl'}
    instructions[1551] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'op': 'load'}
    instructions[1552] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1553] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'op': 'load'}
    instructions[1554] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'op': 'add'}
    instructions[1555] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1556] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'op': 'load'}
    instructions[1557] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'op': 'add'}
    instructions[1558] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'op': 'addl'}
    instructions[1559] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'op': 'load'}
    instructions[1560] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1561] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'op': 'load'}
    instructions[1562] = {5'd17, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'op': 'or'}
    instructions[1563] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'op': 'store'}
    instructions[1564] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'op': 'addl'}
    instructions[1565] = {5'd1, 4'd8, 4'd4, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 4, 'literal': -2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'op': 'addl'}
    instructions[1566] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'op': 'addl'}
    instructions[1567] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'op': 'load'}
    instructions[1568] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'op': 'store'}
    instructions[1569] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'op': 'addl'}
    instructions[1570] = {5'd0, 4'd8, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'op': 'literal'}
    instructions[1571] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'op': 'store'}
    instructions[1572] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'op': 'addl'}
    instructions[1573] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'op': 'addl'}
    instructions[1574] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'op': 'addl'}
    instructions[1575] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'op': 'load'}
    instructions[1576] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1577] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'op': 'load'}
    instructions[1578] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'op': 'add'}
    instructions[1579] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1580] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'op': 'load'}
    instructions[1581] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'op': 'add'}
    instructions[1582] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'op': 'addl'}
    instructions[1583] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1584] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'op': 'load'}
    instructions[1585] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'op': 'store'}
    instructions[1586] = {5'd10, 4'd0, 4'd0, 16'd1587};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413 {'label': 1587, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 413, 'op': 'goto'}
    instructions[1587] = {5'd0, 4'd8, 4'd0, 16'd650};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'literal': 650, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'op': 'literal'}
    instructions[1588] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'op': 'addl'}
    instructions[1589] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'op': 'load'}
    instructions[1590] = {5'd8, 4'd0, 4'd8, 16'd1640};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 8, 'label': 1640, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'op': 'jmp_if_false'}
    instructions[1591] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'op': 'literal'}
    instructions[1592] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'op': 'store'}
    instructions[1593] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'op': 'addl'}
    instructions[1594] = {5'd1, 4'd8, 4'd4, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 4, 'literal': -2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'op': 'addl'}
    instructions[1595] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'op': 'addl'}
    instructions[1596] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'op': 'load'}
    instructions[1597] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'op': 'store'}
    instructions[1598] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'op': 'addl'}
    instructions[1599] = {5'd0, 4'd8, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'op': 'literal'}
    instructions[1600] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'op': 'store'}
    instructions[1601] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'op': 'addl'}
    instructions[1602] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'op': 'addl'}
    instructions[1603] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'op': 'addl'}
    instructions[1604] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'op': 'load'}
    instructions[1605] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1606] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'op': 'load'}
    instructions[1607] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'op': 'add'}
    instructions[1608] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1609] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'op': 'load'}
    instructions[1610] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'op': 'add'}
    instructions[1611] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'op': 'addl'}
    instructions[1612] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'op': 'load'}
    instructions[1613] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1614] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'op': 'load'}
    instructions[1615] = {5'd17, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'op': 'or'}
    instructions[1616] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'op': 'store'}
    instructions[1617] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'op': 'addl'}
    instructions[1618] = {5'd1, 4'd8, 4'd4, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 4, 'literal': -2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'op': 'addl'}
    instructions[1619] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'op': 'addl'}
    instructions[1620] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'op': 'load'}
    instructions[1621] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'op': 'store'}
    instructions[1622] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'op': 'addl'}
    instructions[1623] = {5'd0, 4'd8, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'op': 'literal'}
    instructions[1624] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'op': 'store'}
    instructions[1625] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'op': 'addl'}
    instructions[1626] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'op': 'addl'}
    instructions[1627] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'op': 'addl'}
    instructions[1628] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'op': 'load'}
    instructions[1629] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1630] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'op': 'load'}
    instructions[1631] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'op': 'add'}
    instructions[1632] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1633] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'op': 'load'}
    instructions[1634] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'op': 'add'}
    instructions[1635] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'op': 'addl'}
    instructions[1636] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1637] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'op': 'load'}
    instructions[1638] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'op': 'store'}
    instructions[1639] = {5'd10, 4'd0, 4'd0, 16'd1640};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414 {'label': 1640, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 414, 'op': 'goto'}
    instructions[1640] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 418 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 418, 'op': 'store'}
    instructions[1641] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 418 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 418, 'op': 'addl'}
    instructions[1642] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 418 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 418, 'op': 'store'}
    instructions[1643] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 418 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 418, 'op': 'addl'}
    instructions[1644] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 418 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 418, 'op': 'addl'}
    instructions[1645] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 418 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 418, 'op': 'addl'}
    instructions[1646] = {5'd4, 4'd6, 4'd0, 16'd1952};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 418 {'z': 6, 'label': 1952, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 418, 'op': 'call'}
    instructions[1647] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 418 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 418, 'op': 'addl'}
    instructions[1648] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 418 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 418, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1649] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 418 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 418, 'op': 'load'}
    instructions[1650] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 418 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 418, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1651] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 418 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 418, 'op': 'load'}
    instructions[1652] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 418 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 418, 'op': 'addl'}
    instructions[1653] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 419 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 419, 'op': 'store'}
    instructions[1654] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 419 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 419, 'op': 'addl'}
    instructions[1655] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 419 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 419, 'op': 'store'}
    instructions[1656] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 419 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 419, 'op': 'addl'}
    instructions[1657] = {5'd0, 4'd8, 4'd0, 16'd49320};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 419 {'literal': 49320, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 419, 'op': 'literal'}
    instructions[1658] = {5'd3, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 419 {'a': 8, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 419, 'op': 'literal_hi'}
    instructions[1659] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 419 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 419, 'op': 'store'}
    instructions[1660] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 419 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 419, 'op': 'addl'}
    instructions[1661] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 419 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 419, 'op': 'addl'}
    instructions[1662] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 419 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 419, 'op': 'addl'}
    instructions[1663] = {5'd4, 4'd6, 4'd0, 16'd1962};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 419 {'z': 6, 'label': 1962, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 419, 'op': 'call'}
    instructions[1664] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 419 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 419, 'op': 'addl'}
    instructions[1665] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 419 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 419, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1666] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 419 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 419, 'op': 'load'}
    instructions[1667] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 419 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 419, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1668] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 419 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 419, 'op': 'load'}
    instructions[1669] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 419 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 419, 'op': 'addl'}
    instructions[1670] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 420 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 420, 'op': 'store'}
    instructions[1671] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 420 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 420, 'op': 'addl'}
    instructions[1672] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 420 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 420, 'op': 'store'}
    instructions[1673] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 420 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 420, 'op': 'addl'}
    instructions[1674] = {5'd0, 4'd8, 4'd0, 16'd257};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 420 {'literal': 257, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 420, 'op': 'literal'}
    instructions[1675] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 420 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 420, 'op': 'store'}
    instructions[1676] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 420 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 420, 'op': 'addl'}
    instructions[1677] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 420 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 420, 'op': 'addl'}
    instructions[1678] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 420 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 420, 'op': 'addl'}
    instructions[1679] = {5'd4, 4'd6, 4'd0, 16'd1962};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 420 {'z': 6, 'label': 1962, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 420, 'op': 'call'}
    instructions[1680] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 420 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 420, 'op': 'addl'}
    instructions[1681] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 420 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 420, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1682] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 420 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 420, 'op': 'load'}
    instructions[1683] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 420 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 420, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1684] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 420 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 420, 'op': 'load'}
    instructions[1685] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 420 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 420, 'op': 'addl'}
    instructions[1686] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 421 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 421, 'op': 'store'}
    instructions[1687] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 421 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 421, 'op': 'addl'}
    instructions[1688] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 421 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 421, 'op': 'store'}
    instructions[1689] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 421 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 421, 'op': 'addl'}
    instructions[1690] = {5'd0, 4'd8, 4'd0, 16'd539};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 421 {'literal': 539, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 421, 'op': 'literal'}
    instructions[1691] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 421 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 421, 'op': 'addl'}
    instructions[1692] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 421 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 421, 'op': 'load'}
    instructions[1693] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 421 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 421, 'op': 'store'}
    instructions[1694] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 421 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 421, 'op': 'addl'}
    instructions[1695] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 421 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 421, 'op': 'addl'}
    instructions[1696] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 421 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 421, 'op': 'addl'}
    instructions[1697] = {5'd4, 4'd6, 4'd0, 16'd1962};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 421 {'z': 6, 'label': 1962, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 421, 'op': 'call'}
    instructions[1698] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 421 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 421, 'op': 'addl'}
    instructions[1699] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 421 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 421, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1700] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 421 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 421, 'op': 'load'}
    instructions[1701] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 421 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 421, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1702] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 421 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 421, 'op': 'load'}
    instructions[1703] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 421 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 421, 'op': 'addl'}
    instructions[1704] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 422 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 422, 'op': 'store'}
    instructions[1705] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 422 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 422, 'op': 'addl'}
    instructions[1706] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 422 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 422, 'op': 'store'}
    instructions[1707] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 422 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 422, 'op': 'addl'}
    instructions[1708] = {5'd0, 4'd8, 4'd0, 16'd652};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 422 {'literal': 652, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 422, 'op': 'literal'}
    instructions[1709] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 422 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 422, 'op': 'addl'}
    instructions[1710] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 422 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 422, 'op': 'load'}
    instructions[1711] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 422 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 422, 'op': 'store'}
    instructions[1712] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 422 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 422, 'op': 'addl'}
    instructions[1713] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 422 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 422, 'op': 'addl'}
    instructions[1714] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 422 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 422, 'op': 'addl'}
    instructions[1715] = {5'd4, 4'd6, 4'd0, 16'd1962};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 422 {'z': 6, 'label': 1962, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 422, 'op': 'call'}
    instructions[1716] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 422 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 422, 'op': 'addl'}
    instructions[1717] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 422 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 422, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1718] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 422 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 422, 'op': 'load'}
    instructions[1719] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 422 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 422, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1720] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 422 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 422, 'op': 'load'}
    instructions[1721] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 422 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 422, 'op': 'addl'}
    instructions[1722] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 423 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 423, 'op': 'store'}
    instructions[1723] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 423 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 423, 'op': 'addl'}
    instructions[1724] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 423 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 423, 'op': 'store'}
    instructions[1725] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 423 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 423, 'op': 'addl'}
    instructions[1726] = {5'd0, 4'd8, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 423 {'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 423, 'op': 'literal'}
    instructions[1727] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 423 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 423, 'op': 'store'}
    instructions[1728] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 423 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 423, 'op': 'addl'}
    instructions[1729] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 423 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 423, 'op': 'addl'}
    instructions[1730] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 423 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 423, 'op': 'addl'}
    instructions[1731] = {5'd4, 4'd6, 4'd0, 16'd1962};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 423 {'z': 6, 'label': 1962, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 423, 'op': 'call'}
    instructions[1732] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 423 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 423, 'op': 'addl'}
    instructions[1733] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 423 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 423, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1734] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 423 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 423, 'op': 'load'}
    instructions[1735] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 423 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 423, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1736] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 423 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 423, 'op': 'load'}
    instructions[1737] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 423 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 423, 'op': 'addl'}
    instructions[1738] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424, 'op': 'store'}
    instructions[1739] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424, 'op': 'addl'}
    instructions[1740] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424, 'op': 'store'}
    instructions[1741] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424, 'op': 'addl'}
    instructions[1742] = {5'd0, 4'd8, 4'd0, 16'd20};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424 {'literal': 20, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424, 'op': 'literal'}
    instructions[1743] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424, 'op': 'store'}
    instructions[1744] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424, 'op': 'addl'}
    instructions[1745] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424, 'op': 'addl'}
    instructions[1746] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424, 'op': 'addl'}
    instructions[1747] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424, 'op': 'load'}
    instructions[1748] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1749] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424, 'op': 'load'}
    instructions[1750] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424, 'op': 'add'}
    instructions[1751] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424, 'op': 'store'}
    instructions[1752] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424, 'op': 'addl'}
    instructions[1753] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424, 'op': 'addl'}
    instructions[1754] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424, 'op': 'addl'}
    instructions[1755] = {5'd4, 4'd6, 4'd0, 16'd1962};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424 {'z': 6, 'label': 1962, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424, 'op': 'call'}
    instructions[1756] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424, 'op': 'addl'}
    instructions[1757] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1758] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424, 'op': 'load'}
    instructions[1759] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1760] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424, 'op': 'load'}
    instructions[1761] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 424, 'op': 'addl'}
    instructions[1762] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 426 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 426, 'op': 'literal'}
    instructions[1763] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 426 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 426, 'op': 'store'}
    instructions[1764] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 426 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 426, 'op': 'addl'}
    instructions[1765] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 426 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 426, 'op': 'literal'}
    instructions[1766] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 426 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 426, 'op': 'store'}
    instructions[1767] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 426 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 426, 'op': 'addl'}
    instructions[1768] = {5'd0, 4'd8, 4'd0, 16'd20};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 426 {'literal': 20, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 426, 'op': 'literal'}
    instructions[1769] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 426 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 426, 'op': 'store'}
    instructions[1770] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 426 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 426, 'op': 'addl'}
    instructions[1771] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 426 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 426, 'op': 'addl'}
    instructions[1772] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 426 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 426, 'op': 'addl'}
    instructions[1773] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 426 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 426, 'op': 'load'}
    instructions[1774] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 426 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 426, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1775] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 426 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 426, 'op': 'load'}
    instructions[1776] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 426 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 426, 'op': 'add'}
    instructions[1777] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 426 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 426, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1778] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 426 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 426, 'op': 'load'}
    instructions[1779] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 426 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 426, 'op': 'add'}
    instructions[1780] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 426 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 426, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1781] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 426 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 426, 'op': 'load'}
    instructions[1782] = {5'd18, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 426 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 426, 'op': 'unsigned_shift_right'}
    instructions[1783] = {5'd1, 4'd2, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 426 {'a': 4, 'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 426, 'op': 'addl'}
    instructions[1784] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 426 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 426, 'op': 'store'}
    instructions[1785] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 427 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 427, 'op': 'addl'}
    instructions[1786] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 427 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 427, 'op': 'addl'}
    instructions[1787] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 427 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 427, 'op': 'load'}
    instructions[1788] = {5'd1, 4'd2, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 427 {'a': 4, 'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 427, 'op': 'addl'}
    instructions[1789] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 427 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 427, 'op': 'store'}
    instructions[1790] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428, 'op': 'literal'}
    instructions[1791] = {5'd1, 4'd2, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428 {'a': 4, 'literal': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428, 'op': 'addl'}
    instructions[1792] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428, 'op': 'store'}
    instructions[1793] = {5'd1, 4'd8, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428 {'a': 4, 'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428, 'op': 'addl'}
    instructions[1794] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428, 'op': 'addl'}
    instructions[1795] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428, 'op': 'load'}
    instructions[1796] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428, 'op': 'store'}
    instructions[1797] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428, 'op': 'addl'}
    instructions[1798] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428, 'op': 'addl'}
    instructions[1799] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428, 'op': 'addl'}
    instructions[1800] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428, 'op': 'load'}
    instructions[1801] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1802] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428, 'op': 'load'}
    instructions[1803] = {5'd19, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428, 'op': 'unsigned_greater'}
    instructions[1804] = {5'd8, 4'd0, 4'd8, 16'd1870};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428 {'a': 8, 'label': 1870, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428, 'op': 'jmp_if_false'}
    instructions[1805] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429, 'op': 'store'}
    instructions[1806] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429, 'op': 'addl'}
    instructions[1807] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429, 'op': 'store'}
    instructions[1808] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429, 'op': 'addl'}
    instructions[1809] = {5'd1, 4'd8, 4'd4, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429 {'a': 4, 'literal': -2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429, 'op': 'addl'}
    instructions[1810] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429, 'op': 'addl'}
    instructions[1811] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429, 'op': 'load'}
    instructions[1812] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429, 'op': 'store'}
    instructions[1813] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429, 'op': 'addl'}
    instructions[1814] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429, 'op': 'addl'}
    instructions[1815] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429, 'op': 'addl'}
    instructions[1816] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429, 'op': 'load'}
    instructions[1817] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1818] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429, 'op': 'load'}
    instructions[1819] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429, 'op': 'add'}
    instructions[1820] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429, 'op': 'addl'}
    instructions[1821] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429, 'op': 'load'}
    instructions[1822] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429, 'op': 'store'}
    instructions[1823] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429, 'op': 'addl'}
    instructions[1824] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429, 'op': 'addl'}
    instructions[1825] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429, 'op': 'addl'}
    instructions[1826] = {5'd4, 4'd6, 4'd0, 16'd1962};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429 {'z': 6, 'label': 1962, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429, 'op': 'call'}
    instructions[1827] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429, 'op': 'addl'}
    instructions[1828] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1829] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429, 'op': 'load'}
    instructions[1830] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1831] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429, 'op': 'load'}
    instructions[1832] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 429, 'op': 'addl'}
    instructions[1833] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 430 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 430, 'op': 'addl'}
    instructions[1834] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 430 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 430, 'op': 'addl'}
    instructions[1835] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 430 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 430, 'op': 'load'}
    instructions[1836] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 430 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 430, 'op': 'store'}
    instructions[1837] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 430 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 430, 'op': 'addl'}
    instructions[1838] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 430 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 430, 'op': 'literal'}
    instructions[1839] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 430 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 430, 'op': 'store'}
    instructions[1840] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 430 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 430, 'op': 'addl'}
    instructions[1841] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 430 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 430, 'op': 'addl'}
    instructions[1842] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 430 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 430, 'op': 'addl'}
    instructions[1843] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 430 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 430, 'op': 'load'}
    instructions[1844] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 430 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 430, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1845] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 430 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 430, 'op': 'load'}
    instructions[1846] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 430 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 430, 'op': 'add'}
    instructions[1847] = {5'd1, 4'd2, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 430 {'a': 4, 'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 430, 'op': 'addl'}
    instructions[1848] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 430 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 430, 'op': 'store'}
    instructions[1849] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 430 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 430, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1850] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 430 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 430, 'op': 'load'}
    instructions[1851] = {5'd1, 4'd8, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428 {'a': 4, 'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428, 'op': 'addl'}
    instructions[1852] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428, 'op': 'addl'}
    instructions[1853] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428, 'op': 'load'}
    instructions[1854] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428, 'op': 'store'}
    instructions[1855] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428, 'op': 'addl'}
    instructions[1856] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428, 'op': 'literal'}
    instructions[1857] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428, 'op': 'store'}
    instructions[1858] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428, 'op': 'addl'}
    instructions[1859] = {5'd1, 4'd8, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428 {'a': 4, 'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428, 'op': 'addl'}
    instructions[1860] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428, 'op': 'addl'}
    instructions[1861] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428, 'op': 'load'}
    instructions[1862] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1863] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428, 'op': 'load'}
    instructions[1864] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428, 'op': 'add'}
    instructions[1865] = {5'd1, 4'd2, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428 {'a': 4, 'literal': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428, 'op': 'addl'}
    instructions[1866] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428, 'op': 'store'}
    instructions[1867] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1868] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428, 'op': 'load'}
    instructions[1869] = {5'd10, 4'd0, 4'd0, 16'd1793};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428 {'label': 1793, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 428, 'op': 'goto'}
    instructions[1870] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432, 'op': 'store'}
    instructions[1871] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432, 'op': 'addl'}
    instructions[1872] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432, 'op': 'store'}
    instructions[1873] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432, 'op': 'addl'}
    instructions[1874] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432, 'op': 'addl'}
    instructions[1875] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432, 'op': 'addl'}
    instructions[1876] = {5'd4, 4'd6, 4'd0, 16'd2053};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432 {'z': 6, 'label': 2053, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432, 'op': 'call'}
    instructions[1877] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432, 'op': 'addl'}
    instructions[1878] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1879] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432, 'op': 'load'}
    instructions[1880] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1881] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432, 'op': 'load'}
    instructions[1882] = {5'd0, 4'd2, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432 {'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432, 'op': 'literal'}
    instructions[1883] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432, 'op': 'load'}
    instructions[1884] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432, 'op': 'store'}
    instructions[1885] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432, 'op': 'addl'}
    instructions[1886] = {5'd1, 4'd8, 4'd4, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432 {'a': 4, 'literal': -2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432, 'op': 'addl'}
    instructions[1887] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432, 'op': 'addl'}
    instructions[1888] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432, 'op': 'load'}
    instructions[1889] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432, 'op': 'store'}
    instructions[1890] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432, 'op': 'addl'}
    instructions[1891] = {5'd0, 4'd8, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432 {'literal': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432, 'op': 'literal'}
    instructions[1892] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432, 'op': 'store'}
    instructions[1893] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432, 'op': 'addl'}
    instructions[1894] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432, 'op': 'addl'}
    instructions[1895] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432, 'op': 'addl'}
    instructions[1896] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432, 'op': 'load'}
    instructions[1897] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1898] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432, 'op': 'load'}
    instructions[1899] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432, 'op': 'add'}
    instructions[1900] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1901] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432, 'op': 'load'}
    instructions[1902] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432, 'op': 'add'}
    instructions[1903] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432, 'op': 'addl'}
    instructions[1904] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1905] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432, 'op': 'load'}
    instructions[1906] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 432, 'op': 'store'}
    instructions[1907] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 434 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 434, 'op': 'store'}
    instructions[1908] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 434 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 434, 'op': 'addl'}
    instructions[1909] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 434 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 434, 'op': 'store'}
    instructions[1910] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 434 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 434, 'op': 'addl'}
    instructions[1911] = {5'd1, 4'd8, 4'd4, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 435 {'a': 4, 'literal': -2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 435, 'op': 'addl'}
    instructions[1912] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 435 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 435, 'op': 'addl'}
    instructions[1913] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 435 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 435, 'op': 'load'}
    instructions[1914] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 434 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 434, 'op': 'store'}
    instructions[1915] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 434 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 434, 'op': 'addl'}
    instructions[1916] = {5'd0, 4'd8, 4'd0, 16'd40};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 436 {'literal': 40, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 436, 'op': 'literal'}
    instructions[1917] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 436 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 436, 'op': 'store'}
    instructions[1918] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 436 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 436, 'op': 'addl'}
    instructions[1919] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 436 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 436, 'op': 'addl'}
    instructions[1920] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 436 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 436, 'op': 'addl'}
    instructions[1921] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 436 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 436, 'op': 'load'}
    instructions[1922] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 436 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 436, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1923] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 436 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 436, 'op': 'load'}
    instructions[1924] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 436 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 436, 'op': 'add'}
    instructions[1925] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 434 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 434, 'op': 'store'}
    instructions[1926] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 434 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 434, 'op': 'addl'}
    instructions[1927] = {5'd0, 4'd8, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 437 {'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 437, 'op': 'literal'}
    instructions[1928] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 434 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 434, 'op': 'store'}
    instructions[1929] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 434 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 434, 'op': 'addl'}
    instructions[1930] = {5'd0, 4'd8, 4'd0, 16'd539};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 438 {'literal': 539, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 438, 'op': 'literal'}
    instructions[1931] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 438 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 438, 'op': 'addl'}
    instructions[1932] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 438 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 438, 'op': 'load'}
    instructions[1933] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 434 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 434, 'op': 'store'}
    instructions[1934] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 434 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 434, 'op': 'addl'}
    instructions[1935] = {5'd0, 4'd8, 4'd0, 16'd652};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 439 {'literal': 652, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 439, 'op': 'literal'}
    instructions[1936] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 439 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 439, 'op': 'addl'}
    instructions[1937] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 439 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 439, 'op': 'load'}
    instructions[1938] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 434 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 434, 'op': 'store'}
    instructions[1939] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 434 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 434, 'op': 'addl'}
    instructions[1940] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 434 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 434, 'op': 'addl'}
    instructions[1941] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 434 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 434, 'op': 'addl'}
    instructions[1942] = {5'd4, 4'd6, 4'd0, 16'd2066};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 434 {'z': 6, 'label': 2066, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 434, 'op': 'call'}
    instructions[1943] = {5'd1, 4'd3, 4'd3, -16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 434 {'a': 3, 'literal': -5, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 434, 'op': 'addl'}
    instructions[1944] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 434 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 434, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1945] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 434 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 434, 'op': 'load'}
    instructions[1946] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 434 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 434, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1947] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 434 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 434, 'op': 'load'}
    instructions[1948] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 434 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 434, 'op': 'addl'}
    instructions[1949] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 389 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 389, 'op': 'addl'}
    instructions[1950] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 389 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 389, 'op': 'addl'}
    instructions[1951] = {5'd16, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 389 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 389, 'op': 'return'}
    instructions[1952] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 52 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 52, 'op': 'addl'}
    instructions[1953] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 53 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 53, 'op': 'literal'}
    instructions[1954] = {5'd20, 4'd9, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 53 {'a': 8, 'z': 9, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 53, 'op': 'int_to_long'}
    instructions[1955] = {5'd0, 4'd2, 4'd0, 16'd647};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 53 {'literal': 647, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 53, 'op': 'literal'}
    instructions[1956] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 53 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 53, 'op': 'store'}
    instructions[1957] = {5'd1, 4'd2, 4'd2, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 53 {'a': 2, 'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 53, 'op': 'addl'}
    instructions[1958] = {5'd2, 4'd0, 4'd2, 16'd9};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 53 {'a': 2, 'b': 9, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 53, 'op': 'store'}
    instructions[1959] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 52 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 52, 'op': 'addl'}
    instructions[1960] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 52 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 52, 'op': 'addl'}
    instructions[1961] = {5'd16, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 52 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 52, 'op': 'return'}
    instructions[1962] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 59 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 59, 'op': 'addl'}
    instructions[1963] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 60 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 60, 'op': 'addl'}
    instructions[1964] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 60 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 60, 'op': 'addl'}
    instructions[1965] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 60 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 60, 'op': 'load'}
    instructions[1966] = {5'd0, 4'd9, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 60 {'literal': 0, 'z': 9, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 60, 'op': 'literal'}
    instructions[1967] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 60 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 60, 'op': 'store'}
    instructions[1968] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 60 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 60, 'op': 'addl'}
    instructions[1969] = {5'd2, 4'd0, 4'd3, 16'd9};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 60 {'a': 3, 'comment': 'push', 'b': 9, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 60, 'op': 'store'}
    instructions[1970] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 60 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 60, 'op': 'addl'}
    instructions[1971] = {5'd0, 4'd8, 4'd0, 16'd647};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 60 {'literal': 647, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 60, 'op': 'literal'}
    instructions[1972] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 60 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 60, 'op': 'addl'}
    instructions[1973] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 60 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 60, 'op': 'load'}
    instructions[1974] = {5'd1, 4'd2, 4'd2, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 60 {'a': 2, 'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 60, 'op': 'addl'}
    instructions[1975] = {5'd6, 4'd9, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 60 {'a': 2, 'z': 9, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 60, 'op': 'load'}
    instructions[1976] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 60 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 60, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1977] = {5'd6, 4'd11, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 60 {'a': 3, 'z': 11, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 60, 'op': 'load'}
    instructions[1978] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 60 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 60, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1979] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 60 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 60, 'op': 'load'}
    instructions[1980] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 60 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 60, 'op': 'add'}
    instructions[1981] = {5'd21, 4'd9, 4'd9, 16'd11};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 60 {'a': 9, 'z': 9, 'b': 11, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 60, 'op': 'add_with_carry'}
    instructions[1982] = {5'd0, 4'd2, 4'd0, 16'd647};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 60 {'literal': 647, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 60, 'op': 'literal'}
    instructions[1983] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 60 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 60, 'op': 'store'}
    instructions[1984] = {5'd1, 4'd2, 4'd2, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 60 {'a': 2, 'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 60, 'op': 'addl'}
    instructions[1985] = {5'd2, 4'd0, 4'd2, 16'd9};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 60 {'a': 2, 'b': 9, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 60, 'op': 'store'}
    instructions[1986] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 61 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 61, 'op': 'literal'}
    instructions[1987] = {5'd3, 4'd8, 4'd8, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 61 {'a': 8, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 61, 'op': 'literal_hi'}
    instructions[1988] = {5'd0, 4'd9, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 61 {'literal': 0, 'z': 9, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 61, 'op': 'literal'}
    instructions[1989] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 61 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 61, 'op': 'store'}
    instructions[1990] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 61 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 61, 'op': 'addl'}
    instructions[1991] = {5'd2, 4'd0, 4'd3, 16'd9};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 61 {'a': 3, 'comment': 'push', 'b': 9, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 61, 'op': 'store'}
    instructions[1992] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 61 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 61, 'op': 'addl'}
    instructions[1993] = {5'd0, 4'd8, 4'd0, 16'd647};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 61 {'literal': 647, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 61, 'op': 'literal'}
    instructions[1994] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 61 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 61, 'op': 'addl'}
    instructions[1995] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 61 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 61, 'op': 'load'}
    instructions[1996] = {5'd1, 4'd2, 4'd2, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 61 {'a': 2, 'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 61, 'op': 'addl'}
    instructions[1997] = {5'd6, 4'd9, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 61 {'a': 2, 'z': 9, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 61, 'op': 'load'}
    instructions[1998] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 61 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 61, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1999] = {5'd6, 4'd11, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 61 {'a': 3, 'z': 11, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 61, 'op': 'load'}
    instructions[2000] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 61 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 61, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2001] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 61 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 61, 'op': 'load'}
    instructions[2002] = {5'd22, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 61 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 61, 'op': 'and'}
    instructions[2003] = {5'd22, 4'd9, 4'd9, 16'd11};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 61 {'a': 9, 'z': 9, 'b': 11, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 61, 'op': 'and'}
    instructions[2004] = {5'd17, 4'd8, 4'd8, 16'd9};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 61 {'a': 8, 'z': 8, 'b': 9, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 61, 'op': 'or'}
    instructions[2005] = {5'd8, 4'd0, 4'd8, 16'd2050};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 61 {'a': 8, 'label': 2050, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 61, 'op': 'jmp_if_false'}
    instructions[2006] = {5'd0, 4'd8, 4'd0, 16'd65535};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 62 {'literal': 65535, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 62, 'op': 'literal'}
    instructions[2007] = {5'd3, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 62 {'a': 8, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 62, 'op': 'literal_hi'}
    instructions[2008] = {5'd0, 4'd9, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 62 {'literal': 0, 'z': 9, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 62, 'op': 'literal'}
    instructions[2009] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 62 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 62, 'op': 'store'}
    instructions[2010] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 62 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 62, 'op': 'addl'}
    instructions[2011] = {5'd2, 4'd0, 4'd3, 16'd9};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 62 {'a': 3, 'comment': 'push', 'b': 9, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 62, 'op': 'store'}
    instructions[2012] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 62 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 62, 'op': 'addl'}
    instructions[2013] = {5'd0, 4'd8, 4'd0, 16'd647};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 62 {'literal': 647, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 62, 'op': 'literal'}
    instructions[2014] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 62 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 62, 'op': 'addl'}
    instructions[2015] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 62 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 62, 'op': 'load'}
    instructions[2016] = {5'd1, 4'd2, 4'd2, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 62 {'a': 2, 'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 62, 'op': 'addl'}
    instructions[2017] = {5'd6, 4'd9, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 62 {'a': 2, 'z': 9, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 62, 'op': 'load'}
    instructions[2018] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 62 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 62, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2019] = {5'd6, 4'd11, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 62 {'a': 3, 'z': 11, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 62, 'op': 'load'}
    instructions[2020] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 62 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 62, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2021] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 62 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 62, 'op': 'load'}
    instructions[2022] = {5'd22, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 62 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 62, 'op': 'and'}
    instructions[2023] = {5'd22, 4'd9, 4'd9, 16'd11};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 62 {'a': 9, 'z': 9, 'b': 11, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 62, 'op': 'and'}
    instructions[2024] = {5'd0, 4'd2, 4'd0, 16'd647};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 62 {'literal': 647, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 62, 'op': 'literal'}
    instructions[2025] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 62 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 62, 'op': 'store'}
    instructions[2026] = {5'd1, 4'd2, 4'd2, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 62 {'a': 2, 'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 62, 'op': 'addl'}
    instructions[2027] = {5'd2, 4'd0, 4'd2, 16'd9};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 62 {'a': 2, 'b': 9, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 62, 'op': 'store'}
    instructions[2028] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 63 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 63, 'op': 'literal'}
    instructions[2029] = {5'd0, 4'd9, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 63 {'literal': 0, 'z': 9, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 63, 'op': 'literal'}
    instructions[2030] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 63 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 63, 'op': 'store'}
    instructions[2031] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 63 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 63, 'op': 'addl'}
    instructions[2032] = {5'd2, 4'd0, 4'd3, 16'd9};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 63 {'a': 3, 'comment': 'push', 'b': 9, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 63, 'op': 'store'}
    instructions[2033] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 63 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 63, 'op': 'addl'}
    instructions[2034] = {5'd0, 4'd8, 4'd0, 16'd647};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 63 {'literal': 647, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 63, 'op': 'literal'}
    instructions[2035] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 63 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 63, 'op': 'addl'}
    instructions[2036] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 63 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 63, 'op': 'load'}
    instructions[2037] = {5'd1, 4'd2, 4'd2, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 63 {'a': 2, 'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 63, 'op': 'addl'}
    instructions[2038] = {5'd6, 4'd9, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 63 {'a': 2, 'z': 9, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 63, 'op': 'load'}
    instructions[2039] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 63 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 63, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2040] = {5'd6, 4'd11, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 63 {'a': 3, 'z': 11, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 63, 'op': 'load'}
    instructions[2041] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 63 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 63, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2042] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 63 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 63, 'op': 'load'}
    instructions[2043] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 63 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 63, 'op': 'add'}
    instructions[2044] = {5'd21, 4'd9, 4'd9, 16'd11};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 63 {'a': 9, 'z': 9, 'b': 11, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 63, 'op': 'add_with_carry'}
    instructions[2045] = {5'd0, 4'd2, 4'd0, 16'd647};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 63 {'literal': 647, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 63, 'op': 'literal'}
    instructions[2046] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 63 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 63, 'op': 'store'}
    instructions[2047] = {5'd1, 4'd2, 4'd2, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 63 {'a': 2, 'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 63, 'op': 'addl'}
    instructions[2048] = {5'd2, 4'd0, 4'd2, 16'd9};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 63 {'a': 2, 'b': 9, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 63, 'op': 'store'}
    instructions[2049] = {5'd10, 4'd0, 4'd0, 16'd2050};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 61 {'label': 2050, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 61, 'op': 'goto'}
    instructions[2050] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 59 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 59, 'op': 'addl'}
    instructions[2051] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 59 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 59, 'op': 'addl'}
    instructions[2052] = {5'd16, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 59 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 59, 'op': 'return'}
    instructions[2053] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 70 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 70, 'op': 'addl'}
    instructions[2054] = {5'd0, 4'd8, 4'd0, 16'd647};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 71 {'literal': 647, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 71, 'op': 'literal'}
    instructions[2055] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 71 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 71, 'op': 'addl'}
    instructions[2056] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 71 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 71, 'op': 'load'}
    instructions[2057] = {5'd1, 4'd2, 4'd2, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 71 {'a': 2, 'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 71, 'op': 'addl'}
    instructions[2058] = {5'd6, 4'd9, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 71 {'a': 2, 'z': 9, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 71, 'op': 'load'}
    instructions[2059] = {5'd23, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 71 {'a': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 71, 'op': 'not'}
    instructions[2060] = {5'd23, 4'd9, 4'd9, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 71 {'a': 9, 'z': 9, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 71, 'op': 'not'}
    instructions[2061] = {5'd0, 4'd2, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 71 {'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 71, 'op': 'literal'}
    instructions[2062] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 71 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 71, 'op': 'store'}
    instructions[2063] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 71 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 71, 'op': 'addl'}
    instructions[2064] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 71 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 71, 'op': 'addl'}
    instructions[2065] = {5'd16, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 71 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 71, 'op': 'return'}
    instructions[2066] = {5'd1, 4'd3, 4'd3, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 262 {'a': 3, 'literal': 3, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 262, 'op': 'addl'}
    instructions[2067] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266, 'op': 'store'}
    instructions[2068] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266, 'op': 'addl'}
    instructions[2069] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266, 'op': 'store'}
    instructions[2070] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266, 'op': 'addl'}
    instructions[2071] = {5'd1, 4'd8, 4'd4, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266 {'a': 4, 'literal': -2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266, 'op': 'addl'}
    instructions[2072] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266, 'op': 'addl'}
    instructions[2073] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266, 'op': 'load'}
    instructions[2074] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266, 'op': 'store'}
    instructions[2075] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266, 'op': 'addl'}
    instructions[2076] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266, 'op': 'addl'}
    instructions[2077] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266, 'op': 'addl'}
    instructions[2078] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266, 'op': 'load'}
    instructions[2079] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266, 'op': 'store'}
    instructions[2080] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266, 'op': 'addl'}
    instructions[2081] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266, 'op': 'addl'}
    instructions[2082] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266, 'op': 'addl'}
    instructions[2083] = {5'd4, 4'd6, 4'd0, 16'd2464};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266 {'z': 6, 'label': 2464, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266, 'op': 'call'}
    instructions[2084] = {5'd1, 4'd3, 4'd3, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266 {'a': 3, 'literal': -2, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266, 'op': 'addl'}
    instructions[2085] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2086] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266, 'op': 'load'}
    instructions[2087] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2088] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266, 'op': 'load'}
    instructions[2089] = {5'd0, 4'd2, 4'd0, 16'd589};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266 {'literal': 589, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266, 'op': 'literal'}
    instructions[2090] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266, 'op': 'load'}
    instructions[2091] = {5'd1, 4'd2, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266 {'a': 4, 'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266, 'op': 'addl'}
    instructions[2092] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 266, 'op': 'store'}
    instructions[2093] = {5'd0, 4'd8, 4'd0, 16'd17664};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 269 {'literal': 17664, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 269, 'op': 'literal'}
    instructions[2094] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 269 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 269, 'op': 'store'}
    instructions[2095] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 269 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 269, 'op': 'addl'}
    instructions[2096] = {5'd1, 4'd8, 4'd4, -16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 269 {'a': 4, 'literal': -5, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 269, 'op': 'addl'}
    instructions[2097] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 269 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 269, 'op': 'addl'}
    instructions[2098] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 269 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 269, 'op': 'load'}
    instructions[2099] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 269 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 269, 'op': 'store'}
    instructions[2100] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 269 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 269, 'op': 'addl'}
    instructions[2101] = {5'd0, 4'd8, 4'd0, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 269 {'literal': 7, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 269, 'op': 'literal'}
    instructions[2102] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 269 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 269, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2103] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 269 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 269, 'op': 'load'}
    instructions[2104] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 269 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 269, 'op': 'add'}
    instructions[2105] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 269 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 269, 'op': 'addl'}
    instructions[2106] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 269 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 269, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2107] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 269 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 269, 'op': 'load'}
    instructions[2108] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 269 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 269, 'op': 'store'}
    instructions[2109] = {5'd1, 4'd8, 4'd4, -16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 270 {'a': 4, 'literal': -4, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 270, 'op': 'addl'}
    instructions[2110] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 270 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 270, 'op': 'addl'}
    instructions[2111] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 270 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 270, 'op': 'load'}
    instructions[2112] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 270 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 270, 'op': 'store'}
    instructions[2113] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 270 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 270, 'op': 'addl'}
    instructions[2114] = {5'd1, 4'd8, 4'd4, -16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 270 {'a': 4, 'literal': -5, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 270, 'op': 'addl'}
    instructions[2115] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 270 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 270, 'op': 'addl'}
    instructions[2116] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 270 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 270, 'op': 'load'}
    instructions[2117] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 270 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 270, 'op': 'store'}
    instructions[2118] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 270 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 270, 'op': 'addl'}
    instructions[2119] = {5'd0, 4'd8, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 270 {'literal': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 270, 'op': 'literal'}
    instructions[2120] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 270 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 270, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2121] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 270 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 270, 'op': 'load'}
    instructions[2122] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 270 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 270, 'op': 'add'}
    instructions[2123] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 270 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 270, 'op': 'addl'}
    instructions[2124] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 270 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 270, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2125] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 270 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 270, 'op': 'load'}
    instructions[2126] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 270 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 270, 'op': 'store'}
    instructions[2127] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 271 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 271, 'op': 'literal'}
    instructions[2128] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 271 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 271, 'op': 'store'}
    instructions[2129] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 271 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 271, 'op': 'addl'}
    instructions[2130] = {5'd1, 4'd8, 4'd4, -16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 271 {'a': 4, 'literal': -5, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 271, 'op': 'addl'}
    instructions[2131] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 271 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 271, 'op': 'addl'}
    instructions[2132] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 271 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 271, 'op': 'load'}
    instructions[2133] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 271 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 271, 'op': 'store'}
    instructions[2134] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 271 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 271, 'op': 'addl'}
    instructions[2135] = {5'd0, 4'd8, 4'd0, 16'd9};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 271 {'literal': 9, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 271, 'op': 'literal'}
    instructions[2136] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 271 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 271, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2137] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 271 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 271, 'op': 'load'}
    instructions[2138] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 271 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 271, 'op': 'add'}
    instructions[2139] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 271 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 271, 'op': 'addl'}
    instructions[2140] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 271 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 271, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2141] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 271 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 271, 'op': 'load'}
    instructions[2142] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 271 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 271, 'op': 'store'}
    instructions[2143] = {5'd0, 4'd8, 4'd0, 16'd16384};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 272 {'literal': 16384, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 272, 'op': 'literal'}
    instructions[2144] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 272 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 272, 'op': 'store'}
    instructions[2145] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 272 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 272, 'op': 'addl'}
    instructions[2146] = {5'd1, 4'd8, 4'd4, -16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 272 {'a': 4, 'literal': -5, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 272, 'op': 'addl'}
    instructions[2147] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 272 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 272, 'op': 'addl'}
    instructions[2148] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 272 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 272, 'op': 'load'}
    instructions[2149] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 272 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 272, 'op': 'store'}
    instructions[2150] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 272 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 272, 'op': 'addl'}
    instructions[2151] = {5'd0, 4'd8, 4'd0, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 272 {'literal': 10, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 272, 'op': 'literal'}
    instructions[2152] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 272 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 272, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2153] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 272 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 272, 'op': 'load'}
    instructions[2154] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 272 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 272, 'op': 'add'}
    instructions[2155] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 272 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 272, 'op': 'addl'}
    instructions[2156] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 272 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 272, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2157] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 272 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 272, 'op': 'load'}
    instructions[2158] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 272 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 272, 'op': 'store'}
    instructions[2159] = {5'd1, 4'd8, 4'd4, -16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273 {'a': 4, 'literal': -3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273, 'op': 'addl'}
    instructions[2160] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273, 'op': 'addl'}
    instructions[2161] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273, 'op': 'load'}
    instructions[2162] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273, 'op': 'store'}
    instructions[2163] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273, 'op': 'addl'}
    instructions[2164] = {5'd0, 4'd8, 4'd0, 16'd65280};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273 {'literal': 65280, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273, 'op': 'literal'}
    instructions[2165] = {5'd3, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273 {'a': 8, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273, 'op': 'literal_hi'}
    instructions[2166] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2167] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273, 'op': 'load'}
    instructions[2168] = {5'd17, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273, 'op': 'or'}
    instructions[2169] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273, 'op': 'store'}
    instructions[2170] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273, 'op': 'addl'}
    instructions[2171] = {5'd1, 4'd8, 4'd4, -16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273 {'a': 4, 'literal': -5, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273, 'op': 'addl'}
    instructions[2172] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273, 'op': 'addl'}
    instructions[2173] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273, 'op': 'load'}
    instructions[2174] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273, 'op': 'store'}
    instructions[2175] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273, 'op': 'addl'}
    instructions[2176] = {5'd0, 4'd8, 4'd0, 16'd11};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273 {'literal': 11, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273, 'op': 'literal'}
    instructions[2177] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2178] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273, 'op': 'load'}
    instructions[2179] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273, 'op': 'add'}
    instructions[2180] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273, 'op': 'addl'}
    instructions[2181] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2182] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273, 'op': 'load'}
    instructions[2183] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 273, 'op': 'store'}
    instructions[2184] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 274 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 274, 'op': 'literal'}
    instructions[2185] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 274 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 274, 'op': 'store'}
    instructions[2186] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 274 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 274, 'op': 'addl'}
    instructions[2187] = {5'd1, 4'd8, 4'd4, -16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 274 {'a': 4, 'literal': -5, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 274, 'op': 'addl'}
    instructions[2188] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 274 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 274, 'op': 'addl'}
    instructions[2189] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 274 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 274, 'op': 'load'}
    instructions[2190] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 274 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 274, 'op': 'store'}
    instructions[2191] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 274 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 274, 'op': 'addl'}
    instructions[2192] = {5'd0, 4'd8, 4'd0, 16'd12};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 274 {'literal': 12, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 274, 'op': 'literal'}
    instructions[2193] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 274 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 274, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2194] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 274 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 274, 'op': 'load'}
    instructions[2195] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 274 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 274, 'op': 'add'}
    instructions[2196] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 274 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 274, 'op': 'addl'}
    instructions[2197] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 274 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 274, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2198] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 274 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 274, 'op': 'load'}
    instructions[2199] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 274 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 274, 'op': 'store'}
    instructions[2200] = {5'd0, 4'd8, 4'd0, 16'd49320};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 275 {'literal': 49320, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 275, 'op': 'literal'}
    instructions[2201] = {5'd3, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 275 {'a': 8, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 275, 'op': 'literal_hi'}
    instructions[2202] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 275 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 275, 'op': 'store'}
    instructions[2203] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 275 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 275, 'op': 'addl'}
    instructions[2204] = {5'd1, 4'd8, 4'd4, -16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 275 {'a': 4, 'literal': -5, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 275, 'op': 'addl'}
    instructions[2205] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 275 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 275, 'op': 'addl'}
    instructions[2206] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 275 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 275, 'op': 'load'}
    instructions[2207] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 275 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 275, 'op': 'store'}
    instructions[2208] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 275 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 275, 'op': 'addl'}
    instructions[2209] = {5'd0, 4'd8, 4'd0, 16'd13};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 275 {'literal': 13, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 275, 'op': 'literal'}
    instructions[2210] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 275 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 275, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2211] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 275 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 275, 'op': 'load'}
    instructions[2212] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 275 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 275, 'op': 'add'}
    instructions[2213] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 275 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 275, 'op': 'addl'}
    instructions[2214] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 275 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 275, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2215] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 275 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 275, 'op': 'load'}
    instructions[2216] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 275 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 275, 'op': 'store'}
    instructions[2217] = {5'd0, 4'd8, 4'd0, 16'd257};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 276 {'literal': 257, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 276, 'op': 'literal'}
    instructions[2218] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 276 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 276, 'op': 'store'}
    instructions[2219] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 276 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 276, 'op': 'addl'}
    instructions[2220] = {5'd1, 4'd8, 4'd4, -16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 276 {'a': 4, 'literal': -5, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 276, 'op': 'addl'}
    instructions[2221] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 276 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 276, 'op': 'addl'}
    instructions[2222] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 276 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 276, 'op': 'load'}
    instructions[2223] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 276 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 276, 'op': 'store'}
    instructions[2224] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 276 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 276, 'op': 'addl'}
    instructions[2225] = {5'd0, 4'd8, 4'd0, 16'd14};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 276 {'literal': 14, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 276, 'op': 'literal'}
    instructions[2226] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 276 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 276, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2227] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 276 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 276, 'op': 'load'}
    instructions[2228] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 276 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 276, 'op': 'add'}
    instructions[2229] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 276 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 276, 'op': 'addl'}
    instructions[2230] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 276 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 276, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2231] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 276 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 276, 'op': 'load'}
    instructions[2232] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 276 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 276, 'op': 'store'}
    instructions[2233] = {5'd1, 4'd8, 4'd4, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 277 {'a': 4, 'literal': -2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 277, 'op': 'addl'}
    instructions[2234] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 277 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 277, 'op': 'addl'}
    instructions[2235] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 277 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 277, 'op': 'load'}
    instructions[2236] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 277 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 277, 'op': 'store'}
    instructions[2237] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 277 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 277, 'op': 'addl'}
    instructions[2238] = {5'd1, 4'd8, 4'd4, -16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 277 {'a': 4, 'literal': -5, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 277, 'op': 'addl'}
    instructions[2239] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 277 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 277, 'op': 'addl'}
    instructions[2240] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 277 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 277, 'op': 'load'}
    instructions[2241] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 277 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 277, 'op': 'store'}
    instructions[2242] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 277 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 277, 'op': 'addl'}
    instructions[2243] = {5'd0, 4'd8, 4'd0, 16'd15};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 277 {'literal': 15, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 277, 'op': 'literal'}
    instructions[2244] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 277 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 277, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2245] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 277 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 277, 'op': 'load'}
    instructions[2246] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 277 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 277, 'op': 'add'}
    instructions[2247] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 277 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 277, 'op': 'addl'}
    instructions[2248] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 277 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 277, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2249] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 277 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 277, 'op': 'load'}
    instructions[2250] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 277 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 277, 'op': 'store'}
    instructions[2251] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 278 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 278, 'op': 'addl'}
    instructions[2252] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 278 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 278, 'op': 'addl'}
    instructions[2253] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 278 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 278, 'op': 'load'}
    instructions[2254] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 278 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 278, 'op': 'store'}
    instructions[2255] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 278 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 278, 'op': 'addl'}
    instructions[2256] = {5'd1, 4'd8, 4'd4, -16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 278 {'a': 4, 'literal': -5, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 278, 'op': 'addl'}
    instructions[2257] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 278 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 278, 'op': 'addl'}
    instructions[2258] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 278 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 278, 'op': 'load'}
    instructions[2259] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 278 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 278, 'op': 'store'}
    instructions[2260] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 278 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 278, 'op': 'addl'}
    instructions[2261] = {5'd0, 4'd8, 4'd0, 16'd16};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 278 {'literal': 16, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 278, 'op': 'literal'}
    instructions[2262] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 278 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 278, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2263] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 278 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 278, 'op': 'load'}
    instructions[2264] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 278 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 278, 'op': 'add'}
    instructions[2265] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 278 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 278, 'op': 'addl'}
    instructions[2266] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 278 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 278, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2267] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 278 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 278, 'op': 'load'}
    instructions[2268] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 278 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 278, 'op': 'store'}
    instructions[2269] = {5'd0, 4'd8, 4'd0, 16'd14};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 279 {'literal': 14, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 279, 'op': 'literal'}
    instructions[2270] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 279 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 279, 'op': 'store'}
    instructions[2271] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 279 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 279, 'op': 'addl'}
    instructions[2272] = {5'd1, 4'd8, 4'd4, -16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 279 {'a': 4, 'literal': -4, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 279, 'op': 'addl'}
    instructions[2273] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 279 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 279, 'op': 'addl'}
    instructions[2274] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 279 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 279, 'op': 'load'}
    instructions[2275] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 279 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 279, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2276] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 279 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 279, 'op': 'load'}
    instructions[2277] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 279 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 279, 'op': 'add'}
    instructions[2278] = {5'd1, 4'd2, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 279 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 279, 'op': 'addl'}
    instructions[2279] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 279 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 279, 'op': 'store'}
    instructions[2280] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 282 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 282, 'op': 'store'}
    instructions[2281] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 282 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 282, 'op': 'addl'}
    instructions[2282] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 282 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 282, 'op': 'store'}
    instructions[2283] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 282 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 282, 'op': 'addl'}
    instructions[2284] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 282 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 282, 'op': 'addl'}
    instructions[2285] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 282 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 282, 'op': 'addl'}
    instructions[2286] = {5'd4, 4'd6, 4'd0, 16'd1952};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 282 {'z': 6, 'label': 1952, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 282, 'op': 'call'}
    instructions[2287] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 282 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 282, 'op': 'addl'}
    instructions[2288] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 282 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 282, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2289] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 282 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 282, 'op': 'load'}
    instructions[2290] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 282 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 282, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2291] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 282 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 282, 'op': 'load'}
    instructions[2292] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 282 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 282, 'op': 'addl'}
    instructions[2293] = {5'd0, 4'd8, 4'd0, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283 {'literal': 7, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283, 'op': 'literal'}
    instructions[2294] = {5'd1, 4'd2, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283 {'a': 4, 'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283, 'op': 'addl'}
    instructions[2295] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283, 'op': 'store'}
    instructions[2296] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283, 'op': 'addl'}
    instructions[2297] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283, 'op': 'addl'}
    instructions[2298] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283, 'op': 'load'}
    instructions[2299] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283, 'op': 'store'}
    instructions[2300] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283, 'op': 'addl'}
    instructions[2301] = {5'd0, 4'd8, 4'd0, 16'd16};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283 {'literal': 16, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283, 'op': 'literal'}
    instructions[2302] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2303] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283, 'op': 'load'}
    instructions[2304] = {5'd24, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283, 'op': 'unsigned_greater_equal'}
    instructions[2305] = {5'd8, 4'd0, 4'd8, 16'd2353};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283 {'a': 8, 'label': 2353, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283, 'op': 'jmp_if_false'}
    instructions[2306] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284, 'op': 'store'}
    instructions[2307] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284, 'op': 'addl'}
    instructions[2308] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284, 'op': 'store'}
    instructions[2309] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284, 'op': 'addl'}
    instructions[2310] = {5'd1, 4'd8, 4'd4, -16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284 {'a': 4, 'literal': -5, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284, 'op': 'addl'}
    instructions[2311] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284, 'op': 'addl'}
    instructions[2312] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284, 'op': 'load'}
    instructions[2313] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284, 'op': 'store'}
    instructions[2314] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284, 'op': 'addl'}
    instructions[2315] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284, 'op': 'addl'}
    instructions[2316] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284, 'op': 'addl'}
    instructions[2317] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284, 'op': 'load'}
    instructions[2318] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2319] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284, 'op': 'load'}
    instructions[2320] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284, 'op': 'add'}
    instructions[2321] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284, 'op': 'addl'}
    instructions[2322] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284, 'op': 'load'}
    instructions[2323] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284, 'op': 'store'}
    instructions[2324] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284, 'op': 'addl'}
    instructions[2325] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284, 'op': 'addl'}
    instructions[2326] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284, 'op': 'addl'}
    instructions[2327] = {5'd4, 4'd6, 4'd0, 16'd1962};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284 {'z': 6, 'label': 1962, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284, 'op': 'call'}
    instructions[2328] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284, 'op': 'addl'}
    instructions[2329] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2330] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284, 'op': 'load'}
    instructions[2331] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2332] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284, 'op': 'load'}
    instructions[2333] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 284, 'op': 'addl'}
    instructions[2334] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283, 'op': 'addl'}
    instructions[2335] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283, 'op': 'addl'}
    instructions[2336] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283, 'op': 'load'}
    instructions[2337] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283, 'op': 'store'}
    instructions[2338] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283, 'op': 'addl'}
    instructions[2339] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283, 'op': 'literal'}
    instructions[2340] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283, 'op': 'store'}
    instructions[2341] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283, 'op': 'addl'}
    instructions[2342] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283, 'op': 'addl'}
    instructions[2343] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283, 'op': 'addl'}
    instructions[2344] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283, 'op': 'load'}
    instructions[2345] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2346] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283, 'op': 'load'}
    instructions[2347] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283, 'op': 'add'}
    instructions[2348] = {5'd1, 4'd2, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283 {'a': 4, 'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283, 'op': 'addl'}
    instructions[2349] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283, 'op': 'store'}
    instructions[2350] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2351] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283, 'op': 'load'}
    instructions[2352] = {5'd10, 4'd0, 4'd0, 16'd2296};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283 {'label': 2296, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 283, 'op': 'goto'}
    instructions[2353] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286, 'op': 'store'}
    instructions[2354] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286, 'op': 'addl'}
    instructions[2355] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286, 'op': 'store'}
    instructions[2356] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286, 'op': 'addl'}
    instructions[2357] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286, 'op': 'addl'}
    instructions[2358] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286, 'op': 'addl'}
    instructions[2359] = {5'd4, 4'd6, 4'd0, 16'd2053};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286 {'z': 6, 'label': 2053, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286, 'op': 'call'}
    instructions[2360] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286, 'op': 'addl'}
    instructions[2361] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2362] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286, 'op': 'load'}
    instructions[2363] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2364] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286, 'op': 'load'}
    instructions[2365] = {5'd0, 4'd2, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286 {'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286, 'op': 'literal'}
    instructions[2366] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286, 'op': 'load'}
    instructions[2367] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286, 'op': 'store'}
    instructions[2368] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286, 'op': 'addl'}
    instructions[2369] = {5'd1, 4'd8, 4'd4, -16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286 {'a': 4, 'literal': -5, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286, 'op': 'addl'}
    instructions[2370] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286, 'op': 'addl'}
    instructions[2371] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286, 'op': 'load'}
    instructions[2372] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286, 'op': 'store'}
    instructions[2373] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286, 'op': 'addl'}
    instructions[2374] = {5'd0, 4'd8, 4'd0, 16'd12};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286 {'literal': 12, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286, 'op': 'literal'}
    instructions[2375] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2376] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286, 'op': 'load'}
    instructions[2377] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286, 'op': 'add'}
    instructions[2378] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286, 'op': 'addl'}
    instructions[2379] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2380] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286, 'op': 'load'}
    instructions[2381] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 286, 'op': 'store'}
    instructions[2382] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 289 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 289, 'op': 'addl'}
    instructions[2383] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 289 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 289, 'op': 'addl'}
    instructions[2384] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 289 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 289, 'op': 'load'}
    instructions[2385] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 289 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 289, 'op': 'store'}
    instructions[2386] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 289 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 289, 'op': 'addl'}
    instructions[2387] = {5'd0, 4'd8, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 289 {'literal': 60, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 289, 'op': 'literal'}
    instructions[2388] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 289 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 289, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2389] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 289 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 289, 'op': 'load'}
    instructions[2390] = {5'd19, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 289 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 289, 'op': 'unsigned_greater'}
    instructions[2391] = {5'd8, 4'd0, 4'd8, 16'd2396};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 289 {'a': 8, 'label': 2396, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 289, 'op': 'jmp_if_false'}
    instructions[2392] = {5'd0, 4'd8, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 290 {'literal': 60, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 290, 'op': 'literal'}
    instructions[2393] = {5'd1, 4'd2, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 290 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 290, 'op': 'addl'}
    instructions[2394] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 290 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 290, 'op': 'store'}
    instructions[2395] = {5'd10, 4'd0, 4'd0, 16'd2396};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 289 {'label': 2396, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 289, 'op': 'goto'}
    instructions[2396] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294, 'op': 'store'}
    instructions[2397] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294, 'op': 'addl'}
    instructions[2398] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294, 'op': 'store'}
    instructions[2399] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294, 'op': 'addl'}
    instructions[2400] = {5'd1, 4'd8, 4'd4, -16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 295 {'a': 4, 'literal': -5, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 295, 'op': 'addl'}
    instructions[2401] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 295 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 295, 'op': 'addl'}
    instructions[2402] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 295 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 295, 'op': 'load'}
    instructions[2403] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294, 'op': 'store'}
    instructions[2404] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294, 'op': 'addl'}
    instructions[2405] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 296 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 296, 'op': 'addl'}
    instructions[2406] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 296 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 296, 'op': 'addl'}
    instructions[2407] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 296 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 296, 'op': 'load'}
    instructions[2408] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294, 'op': 'store'}
    instructions[2409] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294, 'op': 'addl'}
    instructions[2410] = {5'd0, 4'd8, 4'd0, 16'd564};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 297 {'literal': 564, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 297, 'op': 'literal'}
    instructions[2411] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 297 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 297, 'op': 'store'}
    instructions[2412] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 297 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 297, 'op': 'addl'}
    instructions[2413] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 297 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 297, 'op': 'addl'}
    instructions[2414] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 297 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 297, 'op': 'addl'}
    instructions[2415] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 297 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 297, 'op': 'load'}
    instructions[2416] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 297 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 297, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2417] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 297 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 297, 'op': 'load'}
    instructions[2418] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 297 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 297, 'op': 'add'}
    instructions[2419] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 297 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 297, 'op': 'addl'}
    instructions[2420] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 297 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 297, 'op': 'load'}
    instructions[2421] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294, 'op': 'store'}
    instructions[2422] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294, 'op': 'addl'}
    instructions[2423] = {5'd0, 4'd8, 4'd0, 16'd592};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 298 {'literal': 592, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 298, 'op': 'literal'}
    instructions[2424] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 298 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 298, 'op': 'store'}
    instructions[2425] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 298 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 298, 'op': 'addl'}
    instructions[2426] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 298 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 298, 'op': 'addl'}
    instructions[2427] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 298 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 298, 'op': 'addl'}
    instructions[2428] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 298 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 298, 'op': 'load'}
    instructions[2429] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 298 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 298, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2430] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 298 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 298, 'op': 'load'}
    instructions[2431] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 298 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 298, 'op': 'add'}
    instructions[2432] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 298 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 298, 'op': 'addl'}
    instructions[2433] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 298 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 298, 'op': 'load'}
    instructions[2434] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294, 'op': 'store'}
    instructions[2435] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294, 'op': 'addl'}
    instructions[2436] = {5'd0, 4'd8, 4'd0, 16'd611};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 299 {'literal': 611, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 299, 'op': 'literal'}
    instructions[2437] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 299 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 299, 'op': 'store'}
    instructions[2438] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 299 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 299, 'op': 'addl'}
    instructions[2439] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 299 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 299, 'op': 'addl'}
    instructions[2440] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 299 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 299, 'op': 'addl'}
    instructions[2441] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 299 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 299, 'op': 'load'}
    instructions[2442] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 299 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 299, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2443] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 299 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 299, 'op': 'load'}
    instructions[2444] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 299 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 299, 'op': 'add'}
    instructions[2445] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 299 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 299, 'op': 'addl'}
    instructions[2446] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 299 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 299, 'op': 'load'}
    instructions[2447] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294, 'op': 'store'}
    instructions[2448] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294, 'op': 'addl'}
    instructions[2449] = {5'd0, 4'd8, 4'd0, 16'd2048};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 300 {'literal': 2048, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 300, 'op': 'literal'}
    instructions[2450] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294, 'op': 'store'}
    instructions[2451] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294, 'op': 'addl'}
    instructions[2452] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294, 'op': 'addl'}
    instructions[2453] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294, 'op': 'addl'}
    instructions[2454] = {5'd4, 4'd6, 4'd0, 16'd3081};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294 {'z': 6, 'label': 3081, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294, 'op': 'call'}
    instructions[2455] = {5'd1, 4'd3, 4'd3, -16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294 {'a': 3, 'literal': -6, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294, 'op': 'addl'}
    instructions[2456] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2457] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294, 'op': 'load'}
    instructions[2458] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2459] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294, 'op': 'load'}
    instructions[2460] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 294, 'op': 'addl'}
    instructions[2461] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 262 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 262, 'op': 'addl'}
    instructions[2462] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 262 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 262, 'op': 'addl'}
    instructions[2463] = {5'd16, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 262 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 262, 'op': 'return'}
    instructions[2464] = {5'd1, 4'd3, 4'd3, 16'd19};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 192 {'a': 3, 'literal': 19, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 192, 'op': 'addl'}
    instructions[2465] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200, 'op': 'literal'}
    instructions[2466] = {5'd1, 4'd2, 4'd4, 16'd18};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200 {'a': 4, 'literal': 18, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200, 'op': 'addl'}
    instructions[2467] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200, 'op': 'store'}
    instructions[2468] = {5'd1, 4'd8, 4'd4, 16'd18};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200 {'a': 4, 'literal': 18, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200, 'op': 'addl'}
    instructions[2469] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200, 'op': 'addl'}
    instructions[2470] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200, 'op': 'load'}
    instructions[2471] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200, 'op': 'store'}
    instructions[2472] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200, 'op': 'addl'}
    instructions[2473] = {5'd0, 4'd8, 4'd0, 16'd16};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200 {'literal': 16, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200, 'op': 'literal'}
    instructions[2474] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2475] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200, 'op': 'load'}
    instructions[2476] = {5'd19, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200, 'op': 'unsigned_greater'}
    instructions[2477] = {5'd8, 4'd0, 4'd8, 16'd2546};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200 {'a': 8, 'label': 2546, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200, 'op': 'jmp_if_false'}
    instructions[2478] = {5'd1, 4'd8, 4'd4, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201 {'a': 4, 'literal': -2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201, 'op': 'addl'}
    instructions[2479] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201, 'op': 'addl'}
    instructions[2480] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201, 'op': 'load'}
    instructions[2481] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201, 'op': 'store'}
    instructions[2482] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201, 'op': 'addl'}
    instructions[2483] = {5'd0, 4'd8, 4'd0, 16'd545};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201 {'literal': 545, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201, 'op': 'literal'}
    instructions[2484] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201, 'op': 'store'}
    instructions[2485] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201, 'op': 'addl'}
    instructions[2486] = {5'd1, 4'd8, 4'd4, 16'd18};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201 {'a': 4, 'literal': 18, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201, 'op': 'addl'}
    instructions[2487] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201, 'op': 'addl'}
    instructions[2488] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201, 'op': 'load'}
    instructions[2489] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2490] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201, 'op': 'load'}
    instructions[2491] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201, 'op': 'add'}
    instructions[2492] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201, 'op': 'addl'}
    instructions[2493] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201, 'op': 'load'}
    instructions[2494] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2495] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201, 'op': 'load'}
    instructions[2496] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201, 'op': 'equal'}
    instructions[2497] = {5'd8, 4'd0, 4'd8, 16'd2517};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201 {'a': 8, 'label': 2517, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201, 'op': 'jmp_if_false'}
    instructions[2498] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201, 'op': 'addl'}
    instructions[2499] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201, 'op': 'addl'}
    instructions[2500] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201, 'op': 'load'}
    instructions[2501] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201, 'op': 'store'}
    instructions[2502] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201, 'op': 'addl'}
    instructions[2503] = {5'd0, 4'd8, 4'd0, 16'd629};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201 {'literal': 629, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201, 'op': 'literal'}
    instructions[2504] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201, 'op': 'store'}
    instructions[2505] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201, 'op': 'addl'}
    instructions[2506] = {5'd1, 4'd8, 4'd4, 16'd18};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201 {'a': 4, 'literal': 18, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201, 'op': 'addl'}
    instructions[2507] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201, 'op': 'addl'}
    instructions[2508] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201, 'op': 'load'}
    instructions[2509] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2510] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201, 'op': 'load'}
    instructions[2511] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201, 'op': 'add'}
    instructions[2512] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201, 'op': 'addl'}
    instructions[2513] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201, 'op': 'load'}
    instructions[2514] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2515] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201, 'op': 'load'}
    instructions[2516] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201, 'op': 'equal'}
    instructions[2517] = {5'd8, 4'd0, 4'd8, 16'd2527};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201 {'a': 8, 'label': 2527, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201, 'op': 'jmp_if_false'}
    instructions[2518] = {5'd1, 4'd8, 4'd4, 16'd18};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 202 {'a': 4, 'literal': 18, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 202, 'op': 'addl'}
    instructions[2519] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 202 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 202, 'op': 'addl'}
    instructions[2520] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 202 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 202, 'op': 'load'}
    instructions[2521] = {5'd0, 4'd2, 4'd0, 16'd589};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 202 {'literal': 589, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 202, 'op': 'literal'}
    instructions[2522] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 202 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 202, 'op': 'store'}
    instructions[2523] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 202 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 202, 'op': 'addl'}
    instructions[2524] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 202 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 202, 'op': 'addl'}
    instructions[2525] = {5'd16, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 202 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 202, 'op': 'return'}
    instructions[2526] = {5'd10, 4'd0, 4'd0, 16'd2527};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201 {'label': 2527, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 201, 'op': 'goto'}
    instructions[2527] = {5'd1, 4'd8, 4'd4, 16'd18};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200 {'a': 4, 'literal': 18, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200, 'op': 'addl'}
    instructions[2528] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200, 'op': 'addl'}
    instructions[2529] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200, 'op': 'load'}
    instructions[2530] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200, 'op': 'store'}
    instructions[2531] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200, 'op': 'addl'}
    instructions[2532] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200, 'op': 'literal'}
    instructions[2533] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200, 'op': 'store'}
    instructions[2534] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200, 'op': 'addl'}
    instructions[2535] = {5'd1, 4'd8, 4'd4, 16'd18};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200 {'a': 4, 'literal': 18, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200, 'op': 'addl'}
    instructions[2536] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200, 'op': 'addl'}
    instructions[2537] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200, 'op': 'load'}
    instructions[2538] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2539] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200, 'op': 'load'}
    instructions[2540] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200, 'op': 'add'}
    instructions[2541] = {5'd1, 4'd2, 4'd4, 16'd18};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200 {'a': 4, 'literal': 18, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200, 'op': 'addl'}
    instructions[2542] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200, 'op': 'store'}
    instructions[2543] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2544] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200, 'op': 'load'}
    instructions[2545] = {5'd10, 4'd0, 4'd0, 16'd2468};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200 {'label': 2468, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 200, 'op': 'goto'}
    instructions[2546] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 207 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 207, 'op': 'literal'}
    instructions[2547] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 207 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 207, 'op': 'store'}
    instructions[2548] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 207 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 207, 'op': 'addl'}
    instructions[2549] = {5'd0, 4'd8, 4'd0, 16'd27};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 207 {'literal': 27, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 207, 'op': 'literal'}
    instructions[2550] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 207 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 207, 'op': 'store'}
    instructions[2551] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 207 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 207, 'op': 'addl'}
    instructions[2552] = {5'd0, 4'd8, 4'd0, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 207 {'literal': 7, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 207, 'op': 'literal'}
    instructions[2553] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 207 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 207, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2554] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 207 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 207, 'op': 'load'}
    instructions[2555] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 207 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 207, 'op': 'add'}
    instructions[2556] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 207 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 207, 'op': 'addl'}
    instructions[2557] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 207 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 207, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2558] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 207 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 207, 'op': 'load'}
    instructions[2559] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 207 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 207, 'op': 'store'}
    instructions[2560] = {5'd0, 4'd8, 4'd0, 16'd2048};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 208 {'literal': 2048, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 208, 'op': 'literal'}
    instructions[2561] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 208 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 208, 'op': 'store'}
    instructions[2562] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 208 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 208, 'op': 'addl'}
    instructions[2563] = {5'd0, 4'd8, 4'd0, 16'd27};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 208 {'literal': 27, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 208, 'op': 'literal'}
    instructions[2564] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 208 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 208, 'op': 'store'}
    instructions[2565] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 208 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 208, 'op': 'addl'}
    instructions[2566] = {5'd0, 4'd8, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 208 {'literal': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 208, 'op': 'literal'}
    instructions[2567] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 208 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 208, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2568] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 208 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 208, 'op': 'load'}
    instructions[2569] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 208 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 208, 'op': 'add'}
    instructions[2570] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 208 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 208, 'op': 'addl'}
    instructions[2571] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 208 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 208, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2572] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 208 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 208, 'op': 'load'}
    instructions[2573] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 208 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 208, 'op': 'store'}
    instructions[2574] = {5'd0, 4'd8, 4'd0, 16'd1540};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 209 {'literal': 1540, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 209, 'op': 'literal'}
    instructions[2575] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 209 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 209, 'op': 'store'}
    instructions[2576] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 209 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 209, 'op': 'addl'}
    instructions[2577] = {5'd0, 4'd8, 4'd0, 16'd27};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 209 {'literal': 27, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 209, 'op': 'literal'}
    instructions[2578] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 209 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 209, 'op': 'store'}
    instructions[2579] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 209 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 209, 'op': 'addl'}
    instructions[2580] = {5'd0, 4'd8, 4'd0, 16'd9};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 209 {'literal': 9, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 209, 'op': 'literal'}
    instructions[2581] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 209 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 209, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2582] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 209 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 209, 'op': 'load'}
    instructions[2583] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 209 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 209, 'op': 'add'}
    instructions[2584] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 209 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 209, 'op': 'addl'}
    instructions[2585] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 209 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 209, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2586] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 209 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 209, 'op': 'load'}
    instructions[2587] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 209 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 209, 'op': 'store'}
    instructions[2588] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 210 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 210, 'op': 'literal'}
    instructions[2589] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 210 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 210, 'op': 'store'}
    instructions[2590] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 210 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 210, 'op': 'addl'}
    instructions[2591] = {5'd0, 4'd8, 4'd0, 16'd27};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 210 {'literal': 27, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 210, 'op': 'literal'}
    instructions[2592] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 210 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 210, 'op': 'store'}
    instructions[2593] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 210 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 210, 'op': 'addl'}
    instructions[2594] = {5'd0, 4'd8, 4'd0, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 210 {'literal': 10, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 210, 'op': 'literal'}
    instructions[2595] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 210 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 210, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2596] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 210 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 210, 'op': 'load'}
    instructions[2597] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 210 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 210, 'op': 'add'}
    instructions[2598] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 210 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 210, 'op': 'addl'}
    instructions[2599] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 210 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 210, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2600] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 210 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 210, 'op': 'load'}
    instructions[2601] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 210 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 210, 'op': 'store'}
    instructions[2602] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 211 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 211, 'op': 'literal'}
    instructions[2603] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 211 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 211, 'op': 'store'}
    instructions[2604] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 211 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 211, 'op': 'addl'}
    instructions[2605] = {5'd0, 4'd8, 4'd0, 16'd27};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 211 {'literal': 27, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 211, 'op': 'literal'}
    instructions[2606] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 211 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 211, 'op': 'store'}
    instructions[2607] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 211 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 211, 'op': 'addl'}
    instructions[2608] = {5'd0, 4'd8, 4'd0, 16'd11};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 211 {'literal': 11, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 211, 'op': 'literal'}
    instructions[2609] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 211 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 211, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2610] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 211 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 211, 'op': 'load'}
    instructions[2611] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 211 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 211, 'op': 'add'}
    instructions[2612] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 211 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 211, 'op': 'addl'}
    instructions[2613] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 211 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 211, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2614] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 211 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 211, 'op': 'load'}
    instructions[2615] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 211 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 211, 'op': 'store'}
    instructions[2616] = {5'd0, 4'd8, 4'd0, 16'd515};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 212 {'literal': 515, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 212, 'op': 'literal'}
    instructions[2617] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 212 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 212, 'op': 'store'}
    instructions[2618] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 212 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 212, 'op': 'addl'}
    instructions[2619] = {5'd0, 4'd8, 4'd0, 16'd27};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 212 {'literal': 27, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 212, 'op': 'literal'}
    instructions[2620] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 212 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 212, 'op': 'store'}
    instructions[2621] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 212 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 212, 'op': 'addl'}
    instructions[2622] = {5'd0, 4'd8, 4'd0, 16'd12};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 212 {'literal': 12, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 212, 'op': 'literal'}
    instructions[2623] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 212 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 212, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2624] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 212 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 212, 'op': 'load'}
    instructions[2625] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 212 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 212, 'op': 'add'}
    instructions[2626] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 212 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 212, 'op': 'addl'}
    instructions[2627] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 212 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 212, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2628] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 212 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 212, 'op': 'load'}
    instructions[2629] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 212 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 212, 'op': 'store'}
    instructions[2630] = {5'd0, 4'd8, 4'd0, 16'd1029};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 213 {'literal': 1029, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 213, 'op': 'literal'}
    instructions[2631] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 213 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 213, 'op': 'store'}
    instructions[2632] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 213 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 213, 'op': 'addl'}
    instructions[2633] = {5'd0, 4'd8, 4'd0, 16'd27};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 213 {'literal': 27, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 213, 'op': 'literal'}
    instructions[2634] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 213 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 213, 'op': 'store'}
    instructions[2635] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 213 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 213, 'op': 'addl'}
    instructions[2636] = {5'd0, 4'd8, 4'd0, 16'd13};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 213 {'literal': 13, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 213, 'op': 'literal'}
    instructions[2637] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 213 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 213, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2638] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 213 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 213, 'op': 'load'}
    instructions[2639] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 213 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 213, 'op': 'add'}
    instructions[2640] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 213 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 213, 'op': 'addl'}
    instructions[2641] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 213 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 213, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2642] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 213 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 213, 'op': 'load'}
    instructions[2643] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 213 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 213, 'op': 'store'}
    instructions[2644] = {5'd0, 4'd8, 4'd0, 16'd49320};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 214 {'literal': 49320, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 214, 'op': 'literal'}
    instructions[2645] = {5'd3, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 214 {'a': 8, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 214, 'op': 'literal_hi'}
    instructions[2646] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 214 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 214, 'op': 'store'}
    instructions[2647] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 214 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 214, 'op': 'addl'}
    instructions[2648] = {5'd0, 4'd8, 4'd0, 16'd27};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 214 {'literal': 27, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 214, 'op': 'literal'}
    instructions[2649] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 214 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 214, 'op': 'store'}
    instructions[2650] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 214 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 214, 'op': 'addl'}
    instructions[2651] = {5'd0, 4'd8, 4'd0, 16'd14};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 214 {'literal': 14, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 214, 'op': 'literal'}
    instructions[2652] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 214 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 214, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2653] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 214 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 214, 'op': 'load'}
    instructions[2654] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 214 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 214, 'op': 'add'}
    instructions[2655] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 214 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 214, 'op': 'addl'}
    instructions[2656] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 214 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 214, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2657] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 214 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 214, 'op': 'load'}
    instructions[2658] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 214 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 214, 'op': 'store'}
    instructions[2659] = {5'd0, 4'd8, 4'd0, 16'd257};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 215 {'literal': 257, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 215, 'op': 'literal'}
    instructions[2660] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 215 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 215, 'op': 'store'}
    instructions[2661] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 215 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 215, 'op': 'addl'}
    instructions[2662] = {5'd0, 4'd8, 4'd0, 16'd27};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 215 {'literal': 27, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 215, 'op': 'literal'}
    instructions[2663] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 215 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 215, 'op': 'store'}
    instructions[2664] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 215 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 215, 'op': 'addl'}
    instructions[2665] = {5'd0, 4'd8, 4'd0, 16'd15};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 215 {'literal': 15, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 215, 'op': 'literal'}
    instructions[2666] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 215 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 215, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2667] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 215 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 215, 'op': 'load'}
    instructions[2668] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 215 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 215, 'op': 'add'}
    instructions[2669] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 215 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 215, 'op': 'addl'}
    instructions[2670] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 215 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 215, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2671] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 215 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 215, 'op': 'load'}
    instructions[2672] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 215 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 215, 'op': 'store'}
    instructions[2673] = {5'd1, 4'd8, 4'd4, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 216 {'a': 4, 'literal': -2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 216, 'op': 'addl'}
    instructions[2674] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 216 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 216, 'op': 'addl'}
    instructions[2675] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 216 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 216, 'op': 'load'}
    instructions[2676] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 216 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 216, 'op': 'store'}
    instructions[2677] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 216 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 216, 'op': 'addl'}
    instructions[2678] = {5'd0, 4'd8, 4'd0, 16'd27};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 216 {'literal': 27, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 216, 'op': 'literal'}
    instructions[2679] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 216 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 216, 'op': 'store'}
    instructions[2680] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 216 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 216, 'op': 'addl'}
    instructions[2681] = {5'd0, 4'd8, 4'd0, 16'd19};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 216 {'literal': 19, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 216, 'op': 'literal'}
    instructions[2682] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 216 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 216, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2683] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 216 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 216, 'op': 'load'}
    instructions[2684] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 216 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 216, 'op': 'add'}
    instructions[2685] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 216 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 216, 'op': 'addl'}
    instructions[2686] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 216 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 216, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2687] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 216 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 216, 'op': 'load'}
    instructions[2688] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 216 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 216, 'op': 'store'}
    instructions[2689] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 217 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 217, 'op': 'addl'}
    instructions[2690] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 217 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 217, 'op': 'addl'}
    instructions[2691] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 217 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 217, 'op': 'load'}
    instructions[2692] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 217 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 217, 'op': 'store'}
    instructions[2693] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 217 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 217, 'op': 'addl'}
    instructions[2694] = {5'd0, 4'd8, 4'd0, 16'd27};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 217 {'literal': 27, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 217, 'op': 'literal'}
    instructions[2695] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 217 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 217, 'op': 'store'}
    instructions[2696] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 217 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 217, 'op': 'addl'}
    instructions[2697] = {5'd0, 4'd8, 4'd0, 16'd20};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 217 {'literal': 20, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 217, 'op': 'literal'}
    instructions[2698] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 217 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 217, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2699] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 217 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 217, 'op': 'load'}
    instructions[2700] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 217 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 217, 'op': 'add'}
    instructions[2701] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 217 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 217, 'op': 'addl'}
    instructions[2702] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 217 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 217, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2703] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 217 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 217, 'op': 'load'}
    instructions[2704] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 217 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 217, 'op': 'store'}
    instructions[2705] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218, 'op': 'store'}
    instructions[2706] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218, 'op': 'addl'}
    instructions[2707] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218, 'op': 'store'}
    instructions[2708] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218, 'op': 'addl'}
    instructions[2709] = {5'd0, 4'd8, 4'd0, 16'd27};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 219 {'literal': 27, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 219, 'op': 'literal'}
    instructions[2710] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218, 'op': 'store'}
    instructions[2711] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218, 'op': 'addl'}
    instructions[2712] = {5'd0, 4'd8, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 220 {'literal': 60, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 220, 'op': 'literal'}
    instructions[2713] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218, 'op': 'store'}
    instructions[2714] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218, 'op': 'addl'}
    instructions[2715] = {5'd0, 4'd8, 4'd0, 16'd65535};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 221 {'literal': 65535, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 221, 'op': 'literal'}
    instructions[2716] = {5'd3, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 221 {'a': 8, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 221, 'op': 'literal_hi'}
    instructions[2717] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218, 'op': 'store'}
    instructions[2718] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218, 'op': 'addl'}
    instructions[2719] = {5'd0, 4'd8, 4'd0, 16'd65535};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 222 {'literal': 65535, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 222, 'op': 'literal'}
    instructions[2720] = {5'd3, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 222 {'a': 8, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 222, 'op': 'literal_hi'}
    instructions[2721] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218, 'op': 'store'}
    instructions[2722] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218, 'op': 'addl'}
    instructions[2723] = {5'd0, 4'd8, 4'd0, 16'd65535};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 223 {'literal': 65535, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 223, 'op': 'literal'}
    instructions[2724] = {5'd3, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 223 {'a': 8, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 223, 'op': 'literal_hi'}
    instructions[2725] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218, 'op': 'store'}
    instructions[2726] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218, 'op': 'addl'}
    instructions[2727] = {5'd0, 4'd8, 4'd0, 16'd2054};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 224 {'literal': 2054, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 224, 'op': 'literal'}
    instructions[2728] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218, 'op': 'store'}
    instructions[2729] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218, 'op': 'addl'}
    instructions[2730] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218, 'op': 'addl'}
    instructions[2731] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218, 'op': 'addl'}
    instructions[2732] = {5'd4, 4'd6, 4'd0, 16'd3081};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218 {'z': 6, 'label': 3081, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218, 'op': 'call'}
    instructions[2733] = {5'd1, 4'd3, 4'd3, -16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218 {'a': 3, 'literal': -6, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218, 'op': 'addl'}
    instructions[2734] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2735] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218, 'op': 'load'}
    instructions[2736] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2737] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218, 'op': 'load'}
    instructions[2738] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 218, 'op': 'addl'}
    instructions[2739] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 229 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 229, 'op': 'store'}
    instructions[2740] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 229 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 229, 'op': 'addl'}
    instructions[2741] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 229 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 229, 'op': 'store'}
    instructions[2742] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 229 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 229, 'op': 'addl'}
    instructions[2743] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 229 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 229, 'op': 'addl'}
    instructions[2744] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 229 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 229, 'op': 'addl'}
    instructions[2745] = {5'd4, 4'd6, 4'd0, 16'd3315};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 229 {'z': 6, 'label': 3315, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 229, 'op': 'call'}
    instructions[2746] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 229 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 229, 'op': 'addl'}
    instructions[2747] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 229 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 229, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2748] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 229 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 229, 'op': 'load'}
    instructions[2749] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 229 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 229, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2750] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 229 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 229, 'op': 'load'}
    instructions[2751] = {5'd0, 4'd2, 4'd0, 16'd540};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 229 {'literal': 540, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 229, 'op': 'literal'}
    instructions[2752] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 229 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 229, 'op': 'load'}
    instructions[2753] = {5'd1, 4'd2, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 229 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 229, 'op': 'addl'}
    instructions[2754] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 229 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 229, 'op': 'store'}
    instructions[2755] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 230 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 230, 'op': 'literal'}
    instructions[2756] = {5'd1, 4'd2, 4'd4, 16'd18};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 230 {'a': 4, 'literal': 18, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 230, 'op': 'addl'}
    instructions[2757] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 230 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 230, 'op': 'store'}
    instructions[2758] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231, 'op': 'literal'}
    instructions[2759] = {5'd1, 4'd2, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231 {'a': 4, 'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231, 'op': 'addl'}
    instructions[2760] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231, 'op': 'store'}
    instructions[2761] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231, 'op': 'addl'}
    instructions[2762] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231, 'op': 'addl'}
    instructions[2763] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231, 'op': 'load'}
    instructions[2764] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231, 'op': 'store'}
    instructions[2765] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231, 'op': 'addl'}
    instructions[2766] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231, 'op': 'addl'}
    instructions[2767] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231, 'op': 'addl'}
    instructions[2768] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231, 'op': 'load'}
    instructions[2769] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2770] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231, 'op': 'load'}
    instructions[2771] = {5'd19, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231, 'op': 'unsigned_greater'}
    instructions[2772] = {5'd8, 4'd0, 4'd8, 16'd2857};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231 {'a': 8, 'label': 2857, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231, 'op': 'jmp_if_false'}
    instructions[2773] = {5'd1, 4'd8, 4'd4, 16'd18};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 233 {'a': 4, 'literal': 18, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 233, 'op': 'addl'}
    instructions[2774] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 233 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 233, 'op': 'addl'}
    instructions[2775] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 233 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 233, 'op': 'load'}
    instructions[2776] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 233 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 233, 'op': 'store'}
    instructions[2777] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 233 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 233, 'op': 'addl'}
    instructions[2778] = {5'd0, 4'd8, 4'd0, 16'd16};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 233 {'literal': 16, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 233, 'op': 'literal'}
    instructions[2779] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 233 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 233, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2780] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 233 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 233, 'op': 'load'}
    instructions[2781] = {5'd19, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 233 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 233, 'op': 'unsigned_greater'}
    instructions[2782] = {5'd8, 4'd0, 4'd8, 16'd2813};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 233 {'a': 8, 'label': 2813, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 233, 'op': 'jmp_if_false'}
    instructions[2783] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234, 'op': 'store'}
    instructions[2784] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234, 'op': 'addl'}
    instructions[2785] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234, 'op': 'store'}
    instructions[2786] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234, 'op': 'addl'}
    instructions[2787] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234, 'op': 'addl'}
    instructions[2788] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234, 'op': 'addl'}
    instructions[2789] = {5'd4, 4'd6, 4'd0, 16'd3315};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234 {'z': 6, 'label': 3315, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234, 'op': 'call'}
    instructions[2790] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234, 'op': 'addl'}
    instructions[2791] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2792] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234, 'op': 'load'}
    instructions[2793] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2794] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234, 'op': 'load'}
    instructions[2795] = {5'd0, 4'd2, 4'd0, 16'd540};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234 {'literal': 540, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234, 'op': 'literal'}
    instructions[2796] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234, 'op': 'load'}
    instructions[2797] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234, 'op': 'store'}
    instructions[2798] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234, 'op': 'addl'}
    instructions[2799] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234, 'op': 'addl'}
    instructions[2800] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234, 'op': 'store'}
    instructions[2801] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234, 'op': 'addl'}
    instructions[2802] = {5'd1, 4'd8, 4'd4, 16'd18};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234 {'a': 4, 'literal': 18, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234, 'op': 'addl'}
    instructions[2803] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234, 'op': 'addl'}
    instructions[2804] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234, 'op': 'load'}
    instructions[2805] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2806] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234, 'op': 'load'}
    instructions[2807] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234, 'op': 'add'}
    instructions[2808] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234, 'op': 'addl'}
    instructions[2809] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2810] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234, 'op': 'load'}
    instructions[2811] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 234, 'op': 'store'}
    instructions[2812] = {5'd10, 4'd0, 4'd0, 16'd2827};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 233 {'label': 2827, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 233, 'op': 'goto'}
    instructions[2813] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 236 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 236, 'op': 'store'}
    instructions[2814] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 236 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 236, 'op': 'addl'}
    instructions[2815] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 236 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 236, 'op': 'store'}
    instructions[2816] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 236 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 236, 'op': 'addl'}
    instructions[2817] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 236 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 236, 'op': 'addl'}
    instructions[2818] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 236 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 236, 'op': 'addl'}
    instructions[2819] = {5'd4, 4'd6, 4'd0, 16'd3315};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 236 {'z': 6, 'label': 3315, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 236, 'op': 'call'}
    instructions[2820] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 236 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 236, 'op': 'addl'}
    instructions[2821] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 236 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 236, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2822] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 236 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 236, 'op': 'load'}
    instructions[2823] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 236 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 236, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2824] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 236 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 236, 'op': 'load'}
    instructions[2825] = {5'd0, 4'd2, 4'd0, 16'd540};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 236 {'literal': 540, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 236, 'op': 'literal'}
    instructions[2826] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 236 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 236, 'op': 'load'}
    instructions[2827] = {5'd1, 4'd8, 4'd4, 16'd18};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 238 {'a': 4, 'literal': 18, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 238, 'op': 'addl'}
    instructions[2828] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 238 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 238, 'op': 'addl'}
    instructions[2829] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 238 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 238, 'op': 'load'}
    instructions[2830] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 238 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 238, 'op': 'store'}
    instructions[2831] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 238 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 238, 'op': 'addl'}
    instructions[2832] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 238 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 238, 'op': 'literal'}
    instructions[2833] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 238 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 238, 'op': 'store'}
    instructions[2834] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 238 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 238, 'op': 'addl'}
    instructions[2835] = {5'd1, 4'd8, 4'd4, 16'd18};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 238 {'a': 4, 'literal': 18, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 238, 'op': 'addl'}
    instructions[2836] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 238 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 238, 'op': 'addl'}
    instructions[2837] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 238 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 238, 'op': 'load'}
    instructions[2838] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 238 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 238, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2839] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 238 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 238, 'op': 'load'}
    instructions[2840] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 238 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 238, 'op': 'add'}
    instructions[2841] = {5'd1, 4'd2, 4'd4, 16'd18};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 238 {'a': 4, 'literal': 18, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 238, 'op': 'addl'}
    instructions[2842] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 238 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 238, 'op': 'store'}
    instructions[2843] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 238 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 238, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2844] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 238 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 238, 'op': 'load'}
    instructions[2845] = {5'd0, 4'd8, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231 {'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231, 'op': 'literal'}
    instructions[2846] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231, 'op': 'store'}
    instructions[2847] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231, 'op': 'addl'}
    instructions[2848] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231, 'op': 'addl'}
    instructions[2849] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231, 'op': 'addl'}
    instructions[2850] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231, 'op': 'load'}
    instructions[2851] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2852] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231, 'op': 'load'}
    instructions[2853] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231, 'op': 'add'}
    instructions[2854] = {5'd1, 4'd2, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231 {'a': 4, 'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231, 'op': 'addl'}
    instructions[2855] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231, 'op': 'store'}
    instructions[2856] = {5'd10, 4'd0, 4'd0, 16'd2761};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231 {'label': 2761, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 231, 'op': 'goto'}
    instructions[2857] = {5'd0, 4'd8, 4'd0, 16'd2054};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242 {'literal': 2054, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242, 'op': 'literal'}
    instructions[2858] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242, 'op': 'store'}
    instructions[2859] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242, 'op': 'addl'}
    instructions[2860] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242, 'op': 'addl'}
    instructions[2861] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242, 'op': 'store'}
    instructions[2862] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242, 'op': 'addl'}
    instructions[2863] = {5'd0, 4'd8, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242 {'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242, 'op': 'literal'}
    instructions[2864] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2865] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242, 'op': 'load'}
    instructions[2866] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242, 'op': 'add'}
    instructions[2867] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242, 'op': 'addl'}
    instructions[2868] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242, 'op': 'load'}
    instructions[2869] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2870] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242, 'op': 'load'}
    instructions[2871] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242, 'op': 'equal'}
    instructions[2872] = {5'd8, 4'd0, 4'd8, 16'd2888};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242 {'a': 8, 'label': 2888, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242, 'op': 'jmp_if_false'}
    instructions[2873] = {5'd0, 4'd8, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242 {'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242, 'op': 'literal'}
    instructions[2874] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242, 'op': 'store'}
    instructions[2875] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242, 'op': 'addl'}
    instructions[2876] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242, 'op': 'addl'}
    instructions[2877] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242, 'op': 'store'}
    instructions[2878] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242, 'op': 'addl'}
    instructions[2879] = {5'd0, 4'd8, 4'd0, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242 {'literal': 10, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242, 'op': 'literal'}
    instructions[2880] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2881] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242, 'op': 'load'}
    instructions[2882] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242, 'op': 'add'}
    instructions[2883] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242, 'op': 'addl'}
    instructions[2884] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242, 'op': 'load'}
    instructions[2885] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2886] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242, 'op': 'load'}
    instructions[2887] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242, 'op': 'equal'}
    instructions[2888] = {5'd8, 4'd0, 4'd8, 16'd3080};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242 {'a': 8, 'label': 3080, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242, 'op': 'jmp_if_false'}
    instructions[2889] = {5'd1, 4'd8, 4'd4, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243 {'a': 4, 'literal': -2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243, 'op': 'addl'}
    instructions[2890] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243, 'op': 'addl'}
    instructions[2891] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243, 'op': 'load'}
    instructions[2892] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243, 'op': 'store'}
    instructions[2893] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243, 'op': 'addl'}
    instructions[2894] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243, 'op': 'addl'}
    instructions[2895] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243, 'op': 'store'}
    instructions[2896] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243, 'op': 'addl'}
    instructions[2897] = {5'd0, 4'd8, 4'd0, 16'd14};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243 {'literal': 14, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243, 'op': 'literal'}
    instructions[2898] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2899] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243, 'op': 'load'}
    instructions[2900] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243, 'op': 'add'}
    instructions[2901] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243, 'op': 'addl'}
    instructions[2902] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243, 'op': 'load'}
    instructions[2903] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2904] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243, 'op': 'load'}
    instructions[2905] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243, 'op': 'equal'}
    instructions[2906] = {5'd8, 4'd0, 4'd8, 16'd2924};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243 {'a': 8, 'label': 2924, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243, 'op': 'jmp_if_false'}
    instructions[2907] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243, 'op': 'addl'}
    instructions[2908] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243, 'op': 'addl'}
    instructions[2909] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243, 'op': 'load'}
    instructions[2910] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243, 'op': 'store'}
    instructions[2911] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243, 'op': 'addl'}
    instructions[2912] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243, 'op': 'addl'}
    instructions[2913] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243, 'op': 'store'}
    instructions[2914] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243, 'op': 'addl'}
    instructions[2915] = {5'd0, 4'd8, 4'd0, 16'd15};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243 {'literal': 15, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243, 'op': 'literal'}
    instructions[2916] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2917] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243, 'op': 'load'}
    instructions[2918] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243, 'op': 'add'}
    instructions[2919] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243, 'op': 'addl'}
    instructions[2920] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243, 'op': 'load'}
    instructions[2921] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2922] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243, 'op': 'load'}
    instructions[2923] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243, 'op': 'equal'}
    instructions[2924] = {5'd8, 4'd0, 4'd8, 16'd3079};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243 {'a': 8, 'label': 3079, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243, 'op': 'jmp_if_false'}
    instructions[2925] = {5'd1, 4'd8, 4'd4, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 244 {'a': 4, 'literal': -2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 244, 'op': 'addl'}
    instructions[2926] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 244 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 244, 'op': 'addl'}
    instructions[2927] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 244 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 244, 'op': 'load'}
    instructions[2928] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 244 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 244, 'op': 'store'}
    instructions[2929] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 244 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 244, 'op': 'addl'}
    instructions[2930] = {5'd0, 4'd8, 4'd0, 16'd545};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 244 {'literal': 545, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 244, 'op': 'literal'}
    instructions[2931] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 244 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 244, 'op': 'store'}
    instructions[2932] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 244 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 244, 'op': 'addl'}
    instructions[2933] = {5'd0, 4'd8, 4'd0, 16'd588};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 244 {'literal': 588, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 244, 'op': 'literal'}
    instructions[2934] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 244 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 244, 'op': 'addl'}
    instructions[2935] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 244 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 244, 'op': 'load'}
    instructions[2936] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 244 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 244, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2937] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 244 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 244, 'op': 'load'}
    instructions[2938] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 244 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 244, 'op': 'add'}
    instructions[2939] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 244 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 244, 'op': 'addl'}
    instructions[2940] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 244 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 244, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2941] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 244 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 244, 'op': 'load'}
    instructions[2942] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 244 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 244, 'op': 'store'}
    instructions[2943] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 245 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 245, 'op': 'addl'}
    instructions[2944] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 245 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 245, 'op': 'addl'}
    instructions[2945] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 245 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 245, 'op': 'load'}
    instructions[2946] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 245 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 245, 'op': 'store'}
    instructions[2947] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 245 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 245, 'op': 'addl'}
    instructions[2948] = {5'd0, 4'd8, 4'd0, 16'd629};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 245 {'literal': 629, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 245, 'op': 'literal'}
    instructions[2949] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 245 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 245, 'op': 'store'}
    instructions[2950] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 245 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 245, 'op': 'addl'}
    instructions[2951] = {5'd0, 4'd8, 4'd0, 16'd588};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 245 {'literal': 588, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 245, 'op': 'literal'}
    instructions[2952] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 245 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 245, 'op': 'addl'}
    instructions[2953] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 245 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 245, 'op': 'load'}
    instructions[2954] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 245 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 245, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2955] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 245 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 245, 'op': 'load'}
    instructions[2956] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 245 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 245, 'op': 'add'}
    instructions[2957] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 245 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 245, 'op': 'addl'}
    instructions[2958] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 245 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 245, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2959] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 245 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 245, 'op': 'load'}
    instructions[2960] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 245 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 245, 'op': 'store'}
    instructions[2961] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246, 'op': 'addl'}
    instructions[2962] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246, 'op': 'store'}
    instructions[2963] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246, 'op': 'addl'}
    instructions[2964] = {5'd0, 4'd8, 4'd0, 16'd11};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246 {'literal': 11, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246, 'op': 'literal'}
    instructions[2965] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2966] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246, 'op': 'load'}
    instructions[2967] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246, 'op': 'add'}
    instructions[2968] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246, 'op': 'addl'}
    instructions[2969] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246, 'op': 'load'}
    instructions[2970] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246, 'op': 'store'}
    instructions[2971] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246, 'op': 'addl'}
    instructions[2972] = {5'd0, 4'd8, 4'd0, 16'd564};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246 {'literal': 564, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246, 'op': 'literal'}
    instructions[2973] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246, 'op': 'store'}
    instructions[2974] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246, 'op': 'addl'}
    instructions[2975] = {5'd0, 4'd8, 4'd0, 16'd588};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246 {'literal': 588, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246, 'op': 'literal'}
    instructions[2976] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246, 'op': 'addl'}
    instructions[2977] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246, 'op': 'load'}
    instructions[2978] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2979] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246, 'op': 'load'}
    instructions[2980] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246, 'op': 'add'}
    instructions[2981] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246, 'op': 'addl'}
    instructions[2982] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2983] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246, 'op': 'load'}
    instructions[2984] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 246, 'op': 'store'}
    instructions[2985] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247, 'op': 'addl'}
    instructions[2986] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247, 'op': 'store'}
    instructions[2987] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247, 'op': 'addl'}
    instructions[2988] = {5'd0, 4'd8, 4'd0, 16'd12};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247 {'literal': 12, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247, 'op': 'literal'}
    instructions[2989] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2990] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247, 'op': 'load'}
    instructions[2991] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247, 'op': 'add'}
    instructions[2992] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247, 'op': 'addl'}
    instructions[2993] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247, 'op': 'load'}
    instructions[2994] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247, 'op': 'store'}
    instructions[2995] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247, 'op': 'addl'}
    instructions[2996] = {5'd0, 4'd8, 4'd0, 16'd592};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247 {'literal': 592, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247, 'op': 'literal'}
    instructions[2997] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247, 'op': 'store'}
    instructions[2998] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247, 'op': 'addl'}
    instructions[2999] = {5'd0, 4'd8, 4'd0, 16'd588};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247 {'literal': 588, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247, 'op': 'literal'}
    instructions[3000] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247, 'op': 'addl'}
    instructions[3001] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247, 'op': 'load'}
    instructions[3002] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3003] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247, 'op': 'load'}
    instructions[3004] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247, 'op': 'add'}
    instructions[3005] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247, 'op': 'addl'}
    instructions[3006] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3007] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247, 'op': 'load'}
    instructions[3008] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 247, 'op': 'store'}
    instructions[3009] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248, 'op': 'addl'}
    instructions[3010] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248, 'op': 'store'}
    instructions[3011] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248, 'op': 'addl'}
    instructions[3012] = {5'd0, 4'd8, 4'd0, 16'd13};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248 {'literal': 13, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248, 'op': 'literal'}
    instructions[3013] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3014] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248, 'op': 'load'}
    instructions[3015] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248, 'op': 'add'}
    instructions[3016] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248, 'op': 'addl'}
    instructions[3017] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248, 'op': 'load'}
    instructions[3018] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248, 'op': 'store'}
    instructions[3019] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248, 'op': 'addl'}
    instructions[3020] = {5'd0, 4'd8, 4'd0, 16'd611};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248 {'literal': 611, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248, 'op': 'literal'}
    instructions[3021] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248, 'op': 'store'}
    instructions[3022] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248, 'op': 'addl'}
    instructions[3023] = {5'd0, 4'd8, 4'd0, 16'd588};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248 {'literal': 588, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248, 'op': 'literal'}
    instructions[3024] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248, 'op': 'addl'}
    instructions[3025] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248, 'op': 'load'}
    instructions[3026] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3027] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248, 'op': 'load'}
    instructions[3028] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248, 'op': 'add'}
    instructions[3029] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248, 'op': 'addl'}
    instructions[3030] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3031] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248, 'op': 'load'}
    instructions[3032] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 248, 'op': 'store'}
    instructions[3033] = {5'd0, 4'd8, 4'd0, 16'd588};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 249 {'literal': 588, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 249, 'op': 'literal'}
    instructions[3034] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 249 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 249, 'op': 'addl'}
    instructions[3035] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 249 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 249, 'op': 'load'}
    instructions[3036] = {5'd1, 4'd2, 4'd4, 16'd18};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 249 {'a': 4, 'literal': 18, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 249, 'op': 'addl'}
    instructions[3037] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 249 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 249, 'op': 'store'}
    instructions[3038] = {5'd0, 4'd8, 4'd0, 16'd588};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 250 {'literal': 588, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 250, 'op': 'literal'}
    instructions[3039] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 250 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 250, 'op': 'addl'}
    instructions[3040] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 250 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 250, 'op': 'load'}
    instructions[3041] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 250 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 250, 'op': 'store'}
    instructions[3042] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 250 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 250, 'op': 'addl'}
    instructions[3043] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 250 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 250, 'op': 'literal'}
    instructions[3044] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 250 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 250, 'op': 'store'}
    instructions[3045] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 250 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 250, 'op': 'addl'}
    instructions[3046] = {5'd0, 4'd8, 4'd0, 16'd588};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 250 {'literal': 588, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 250, 'op': 'literal'}
    instructions[3047] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 250 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 250, 'op': 'addl'}
    instructions[3048] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 250 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 250, 'op': 'load'}
    instructions[3049] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 250 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 250, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3050] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 250 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 250, 'op': 'load'}
    instructions[3051] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 250 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 250, 'op': 'add'}
    instructions[3052] = {5'd0, 4'd2, 4'd0, 16'd588};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 250 {'literal': 588, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 250, 'op': 'literal'}
    instructions[3053] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 250 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 250, 'op': 'store'}
    instructions[3054] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 250 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 250, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3055] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 250 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 250, 'op': 'load'}
    instructions[3056] = {5'd0, 4'd8, 4'd0, 16'd16};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 251 {'literal': 16, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 251, 'op': 'literal'}
    instructions[3057] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 251 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 251, 'op': 'store'}
    instructions[3058] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 251 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 251, 'op': 'addl'}
    instructions[3059] = {5'd0, 4'd8, 4'd0, 16'd588};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 251 {'literal': 588, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 251, 'op': 'literal'}
    instructions[3060] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 251 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 251, 'op': 'addl'}
    instructions[3061] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 251 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 251, 'op': 'load'}
    instructions[3062] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 251 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 251, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3063] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 251 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 251, 'op': 'load'}
    instructions[3064] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 251 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 251, 'op': 'equal'}
    instructions[3065] = {5'd8, 4'd0, 4'd8, 16'd3070};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 251 {'a': 8, 'label': 3070, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 251, 'op': 'jmp_if_false'}
    instructions[3066] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 251 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 251, 'op': 'literal'}
    instructions[3067] = {5'd0, 4'd2, 4'd0, 16'd588};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 251 {'literal': 588, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 251, 'op': 'literal'}
    instructions[3068] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 251 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 251, 'op': 'store'}
    instructions[3069] = {5'd10, 4'd0, 4'd0, 16'd3070};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 251 {'label': 3070, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 251, 'op': 'goto'}
    instructions[3070] = {5'd1, 4'd8, 4'd4, 16'd18};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 252 {'a': 4, 'literal': 18, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 252, 'op': 'addl'}
    instructions[3071] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 252 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 252, 'op': 'addl'}
    instructions[3072] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 252 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 252, 'op': 'load'}
    instructions[3073] = {5'd0, 4'd2, 4'd0, 16'd589};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 252 {'literal': 589, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 252, 'op': 'literal'}
    instructions[3074] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 252 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 252, 'op': 'store'}
    instructions[3075] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 252 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 252, 'op': 'addl'}
    instructions[3076] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 252 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 252, 'op': 'addl'}
    instructions[3077] = {5'd16, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 252 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 252, 'op': 'return'}
    instructions[3078] = {5'd10, 4'd0, 4'd0, 16'd3079};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243 {'label': 3079, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 243, 'op': 'goto'}
    instructions[3079] = {5'd10, 4'd0, 4'd0, 16'd3080};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242 {'label': 3080, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 242, 'op': 'goto'}
    instructions[3080] = {5'd10, 4'd0, 4'd0, 16'd2739};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 227 {'label': 2739, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 227, 'op': 'goto'}
    instructions[3081] = {5'd1, 4'd3, 4'd3, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 102 {'a': 3, 'literal': 2, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 102, 'op': 'addl'}
    instructions[3082] = {5'd1, 4'd8, 4'd4, -16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 113 {'a': 4, 'literal': -4, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 113, 'op': 'addl'}
    instructions[3083] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 113 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 113, 'op': 'addl'}
    instructions[3084] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 113 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 113, 'op': 'load'}
    instructions[3085] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 113 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 113, 'op': 'store'}
    instructions[3086] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 113 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 113, 'op': 'addl'}
    instructions[3087] = {5'd1, 4'd8, 4'd4, -16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 113 {'a': 4, 'literal': -6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 113, 'op': 'addl'}
    instructions[3088] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 113 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 113, 'op': 'addl'}
    instructions[3089] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 113 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 113, 'op': 'load'}
    instructions[3090] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 113 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 113, 'op': 'store'}
    instructions[3091] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 113 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 113, 'op': 'addl'}
    instructions[3092] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 113 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 113, 'op': 'literal'}
    instructions[3093] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 113 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 113, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3094] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 113 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 113, 'op': 'load'}
    instructions[3095] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 113 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 113, 'op': 'add'}
    instructions[3096] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 113 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 113, 'op': 'addl'}
    instructions[3097] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 113 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 113, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3098] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 113 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 113, 'op': 'load'}
    instructions[3099] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 113 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 113, 'op': 'store'}
    instructions[3100] = {5'd1, 4'd8, 4'd4, -16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 114 {'a': 4, 'literal': -3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 114, 'op': 'addl'}
    instructions[3101] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 114 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 114, 'op': 'addl'}
    instructions[3102] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 114 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 114, 'op': 'load'}
    instructions[3103] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 114 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 114, 'op': 'store'}
    instructions[3104] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 114 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 114, 'op': 'addl'}
    instructions[3105] = {5'd1, 4'd8, 4'd4, -16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 114 {'a': 4, 'literal': -6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 114, 'op': 'addl'}
    instructions[3106] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 114 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 114, 'op': 'addl'}
    instructions[3107] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 114 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 114, 'op': 'load'}
    instructions[3108] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 114 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 114, 'op': 'store'}
    instructions[3109] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 114 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 114, 'op': 'addl'}
    instructions[3110] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 114 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 114, 'op': 'literal'}
    instructions[3111] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 114 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 114, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3112] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 114 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 114, 'op': 'load'}
    instructions[3113] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 114 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 114, 'op': 'add'}
    instructions[3114] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 114 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 114, 'op': 'addl'}
    instructions[3115] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 114 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 114, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3116] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 114 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 114, 'op': 'load'}
    instructions[3117] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 114 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 114, 'op': 'store'}
    instructions[3118] = {5'd1, 4'd8, 4'd4, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 115 {'a': 4, 'literal': -2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 115, 'op': 'addl'}
    instructions[3119] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 115 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 115, 'op': 'addl'}
    instructions[3120] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 115 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 115, 'op': 'load'}
    instructions[3121] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 115 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 115, 'op': 'store'}
    instructions[3122] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 115 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 115, 'op': 'addl'}
    instructions[3123] = {5'd1, 4'd8, 4'd4, -16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 115 {'a': 4, 'literal': -6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 115, 'op': 'addl'}
    instructions[3124] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 115 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 115, 'op': 'addl'}
    instructions[3125] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 115 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 115, 'op': 'load'}
    instructions[3126] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 115 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 115, 'op': 'store'}
    instructions[3127] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 115 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 115, 'op': 'addl'}
    instructions[3128] = {5'd0, 4'd8, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 115 {'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 115, 'op': 'literal'}
    instructions[3129] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 115 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 115, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3130] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 115 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 115, 'op': 'load'}
    instructions[3131] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 115 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 115, 'op': 'add'}
    instructions[3132] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 115 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 115, 'op': 'addl'}
    instructions[3133] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 115 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 115, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3134] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 115 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 115, 'op': 'load'}
    instructions[3135] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 115 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 115, 'op': 'store'}
    instructions[3136] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 116 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 116, 'op': 'literal'}
    instructions[3137] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 116 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 116, 'op': 'store'}
    instructions[3138] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 116 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 116, 'op': 'addl'}
    instructions[3139] = {5'd1, 4'd8, 4'd4, -16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 116 {'a': 4, 'literal': -6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 116, 'op': 'addl'}
    instructions[3140] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 116 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 116, 'op': 'addl'}
    instructions[3141] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 116 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 116, 'op': 'load'}
    instructions[3142] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 116 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 116, 'op': 'store'}
    instructions[3143] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 116 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 116, 'op': 'addl'}
    instructions[3144] = {5'd0, 4'd8, 4'd0, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 116 {'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 116, 'op': 'literal'}
    instructions[3145] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 116 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 116, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3146] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 116 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 116, 'op': 'load'}
    instructions[3147] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 116 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 116, 'op': 'add'}
    instructions[3148] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 116 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 116, 'op': 'addl'}
    instructions[3149] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 116 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 116, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3150] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 116 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 116, 'op': 'load'}
    instructions[3151] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 116 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 116, 'op': 'store'}
    instructions[3152] = {5'd0, 4'd8, 4'd0, 16'd515};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 117 {'literal': 515, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 117, 'op': 'literal'}
    instructions[3153] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 117 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 117, 'op': 'store'}
    instructions[3154] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 117 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 117, 'op': 'addl'}
    instructions[3155] = {5'd1, 4'd8, 4'd4, -16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 117 {'a': 4, 'literal': -6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 117, 'op': 'addl'}
    instructions[3156] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 117 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 117, 'op': 'addl'}
    instructions[3157] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 117 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 117, 'op': 'load'}
    instructions[3158] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 117 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 117, 'op': 'store'}
    instructions[3159] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 117 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 117, 'op': 'addl'}
    instructions[3160] = {5'd0, 4'd8, 4'd0, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 117 {'literal': 4, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 117, 'op': 'literal'}
    instructions[3161] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 117 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 117, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3162] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 117 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 117, 'op': 'load'}
    instructions[3163] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 117 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 117, 'op': 'add'}
    instructions[3164] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 117 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 117, 'op': 'addl'}
    instructions[3165] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 117 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 117, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3166] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 117 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 117, 'op': 'load'}
    instructions[3167] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 117 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 117, 'op': 'store'}
    instructions[3168] = {5'd0, 4'd8, 4'd0, 16'd1029};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 118 {'literal': 1029, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 118, 'op': 'literal'}
    instructions[3169] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 118 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 118, 'op': 'store'}
    instructions[3170] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 118 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 118, 'op': 'addl'}
    instructions[3171] = {5'd1, 4'd8, 4'd4, -16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 118 {'a': 4, 'literal': -6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 118, 'op': 'addl'}
    instructions[3172] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 118 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 118, 'op': 'addl'}
    instructions[3173] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 118 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 118, 'op': 'load'}
    instructions[3174] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 118 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 118, 'op': 'store'}
    instructions[3175] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 118 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 118, 'op': 'addl'}
    instructions[3176] = {5'd0, 4'd8, 4'd0, 16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 118 {'literal': 5, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 118, 'op': 'literal'}
    instructions[3177] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 118 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 118, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3178] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 118 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 118, 'op': 'load'}
    instructions[3179] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 118 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 118, 'op': 'add'}
    instructions[3180] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 118 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 118, 'op': 'addl'}
    instructions[3181] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 118 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 118, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3182] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 118 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 118, 'op': 'load'}
    instructions[3183] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 118 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 118, 'op': 'store'}
    instructions[3184] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 119 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 119, 'op': 'addl'}
    instructions[3185] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 119 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 119, 'op': 'addl'}
    instructions[3186] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 119 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 119, 'op': 'load'}
    instructions[3187] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 119 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 119, 'op': 'store'}
    instructions[3188] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 119 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 119, 'op': 'addl'}
    instructions[3189] = {5'd1, 4'd8, 4'd4, -16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 119 {'a': 4, 'literal': -6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 119, 'op': 'addl'}
    instructions[3190] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 119 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 119, 'op': 'addl'}
    instructions[3191] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 119 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 119, 'op': 'load'}
    instructions[3192] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 119 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 119, 'op': 'store'}
    instructions[3193] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 119 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 119, 'op': 'addl'}
    instructions[3194] = {5'd0, 4'd8, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 119 {'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 119, 'op': 'literal'}
    instructions[3195] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 119 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 119, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3196] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 119 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 119, 'op': 'load'}
    instructions[3197] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 119 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 119, 'op': 'add'}
    instructions[3198] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 119 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 119, 'op': 'addl'}
    instructions[3199] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 119 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 119, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3200] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 119 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 119, 'op': 'load'}
    instructions[3201] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 119 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 119, 'op': 'store'}
    instructions[3202] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 121 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 121, 'op': 'store'}
    instructions[3203] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 121 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 121, 'op': 'addl'}
    instructions[3204] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 121 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 121, 'op': 'store'}
    instructions[3205] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 121 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 121, 'op': 'addl'}
    instructions[3206] = {5'd1, 4'd8, 4'd4, -16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 121 {'a': 4, 'literal': -5, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 121, 'op': 'addl'}
    instructions[3207] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 121 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 121, 'op': 'addl'}
    instructions[3208] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 121 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 121, 'op': 'load'}
    instructions[3209] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 121 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 121, 'op': 'store'}
    instructions[3210] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 121 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 121, 'op': 'addl'}
    instructions[3211] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 121 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 121, 'op': 'addl'}
    instructions[3212] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 121 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 121, 'op': 'addl'}
    instructions[3213] = {5'd4, 4'd6, 4'd0, 16'd3299};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 121 {'z': 6, 'label': 3299, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 121, 'op': 'call'}
    instructions[3214] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 121 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 121, 'op': 'addl'}
    instructions[3215] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 121 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 121, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3216] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 121 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 121, 'op': 'load'}
    instructions[3217] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 121 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 121, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3218] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 121 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 121, 'op': 'load'}
    instructions[3219] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 121 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 121, 'op': 'addl'}
    instructions[3220] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 122 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 122, 'op': 'literal'}
    instructions[3221] = {5'd1, 4'd2, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 122 {'a': 4, 'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 122, 'op': 'addl'}
    instructions[3222] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 122 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 122, 'op': 'store'}
    instructions[3223] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123, 'op': 'literal'}
    instructions[3224] = {5'd1, 4'd2, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123, 'op': 'addl'}
    instructions[3225] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123, 'op': 'store'}
    instructions[3226] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123, 'op': 'addl'}
    instructions[3227] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123, 'op': 'addl'}
    instructions[3228] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123, 'op': 'load'}
    instructions[3229] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123, 'op': 'store'}
    instructions[3230] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123, 'op': 'addl'}
    instructions[3231] = {5'd1, 4'd8, 4'd4, -16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123 {'a': 4, 'literal': -5, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123, 'op': 'addl'}
    instructions[3232] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123, 'op': 'addl'}
    instructions[3233] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123, 'op': 'load'}
    instructions[3234] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3235] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123, 'op': 'load'}
    instructions[3236] = {5'd19, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123, 'op': 'unsigned_greater'}
    instructions[3237] = {5'd8, 4'd0, 4'd8, 16'd3296};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123 {'a': 8, 'label': 3296, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123, 'op': 'jmp_if_false'}
    instructions[3238] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124, 'op': 'store'}
    instructions[3239] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124, 'op': 'addl'}
    instructions[3240] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124, 'op': 'store'}
    instructions[3241] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124, 'op': 'addl'}
    instructions[3242] = {5'd1, 4'd8, 4'd4, -16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124 {'a': 4, 'literal': -6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124, 'op': 'addl'}
    instructions[3243] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124, 'op': 'addl'}
    instructions[3244] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124, 'op': 'load'}
    instructions[3245] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124, 'op': 'store'}
    instructions[3246] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124, 'op': 'addl'}
    instructions[3247] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124, 'op': 'addl'}
    instructions[3248] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124, 'op': 'addl'}
    instructions[3249] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124, 'op': 'load'}
    instructions[3250] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3251] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124, 'op': 'load'}
    instructions[3252] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124, 'op': 'add'}
    instructions[3253] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124, 'op': 'addl'}
    instructions[3254] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124, 'op': 'load'}
    instructions[3255] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124, 'op': 'store'}
    instructions[3256] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124, 'op': 'addl'}
    instructions[3257] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124, 'op': 'addl'}
    instructions[3258] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124, 'op': 'addl'}
    instructions[3259] = {5'd4, 4'd6, 4'd0, 16'd3299};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124 {'z': 6, 'label': 3299, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124, 'op': 'call'}
    instructions[3260] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124, 'op': 'addl'}
    instructions[3261] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3262] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124, 'op': 'load'}
    instructions[3263] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3264] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124, 'op': 'load'}
    instructions[3265] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 124, 'op': 'addl'}
    instructions[3266] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 125 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 125, 'op': 'addl'}
    instructions[3267] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 125 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 125, 'op': 'addl'}
    instructions[3268] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 125 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 125, 'op': 'load'}
    instructions[3269] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 125 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 125, 'op': 'store'}
    instructions[3270] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 125 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 125, 'op': 'addl'}
    instructions[3271] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 125 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 125, 'op': 'literal'}
    instructions[3272] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 125 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 125, 'op': 'store'}
    instructions[3273] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 125 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 125, 'op': 'addl'}
    instructions[3274] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 125 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 125, 'op': 'addl'}
    instructions[3275] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 125 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 125, 'op': 'addl'}
    instructions[3276] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 125 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 125, 'op': 'load'}
    instructions[3277] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 125 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 125, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3278] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 125 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 125, 'op': 'load'}
    instructions[3279] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 125 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 125, 'op': 'add'}
    instructions[3280] = {5'd1, 4'd2, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 125 {'a': 4, 'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 125, 'op': 'addl'}
    instructions[3281] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 125 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 125, 'op': 'store'}
    instructions[3282] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 125 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 125, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3283] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 125 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 125, 'op': 'load'}
    instructions[3284] = {5'd0, 4'd8, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123 {'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123, 'op': 'literal'}
    instructions[3285] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123, 'op': 'store'}
    instructions[3286] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123, 'op': 'addl'}
    instructions[3287] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123, 'op': 'addl'}
    instructions[3288] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123, 'op': 'addl'}
    instructions[3289] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123, 'op': 'load'}
    instructions[3290] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3291] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123, 'op': 'load'}
    instructions[3292] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123, 'op': 'add'}
    instructions[3293] = {5'd1, 4'd2, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123, 'op': 'addl'}
    instructions[3294] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123, 'op': 'store'}
    instructions[3295] = {5'd10, 4'd0, 4'd0, 16'd3226};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123 {'label': 3226, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 123, 'op': 'goto'}
    instructions[3296] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 102 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 102, 'op': 'addl'}
    instructions[3297] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 102 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 102, 'op': 'addl'}
    instructions[3298] = {5'd16, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 102 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 102, 'op': 'return'}
    instructions[3299] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 18 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 18, 'op': 'addl'}
    instructions[3300] = {5'd0, 4'd8, 4'd0, 16'd585};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 19 {'literal': 585, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 19, 'op': 'literal'}
    instructions[3301] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 19 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 19, 'op': 'addl'}
    instructions[3302] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 19 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 19, 'op': 'load'}
    instructions[3303] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 19 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 19, 'op': 'store'}
    instructions[3304] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 19 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 19, 'op': 'addl'}
    instructions[3305] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 19 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 19, 'op': 'addl'}
    instructions[3306] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 19 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 19, 'op': 'addl'}
    instructions[3307] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 19 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 19, 'op': 'load'}
    instructions[3308] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 19 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 19, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3309] = {5'd6, 4'd0, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 19 {'a': 3, 'z': 0, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 19, 'op': 'load'}
    instructions[3310] = {5'd25, 4'd0, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 19 {'a': 0, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 19, 'op': 'write'}
    instructions[3311] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 19 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 19, 'op': 'addl'}
    instructions[3312] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 18 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 18, 'op': 'addl'}
    instructions[3313] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 18 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 18, 'op': 'addl'}
    instructions[3314] = {5'd16, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 18 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 18, 'op': 'return'}
    instructions[3315] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 24 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 24, 'op': 'addl'}
    instructions[3316] = {5'd0, 4'd8, 4'd0, 16'd654};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 25 {'literal': 654, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 25, 'op': 'literal'}
    instructions[3317] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 25 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 25, 'op': 'addl'}
    instructions[3318] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 25 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 25, 'op': 'load'}
    instructions[3319] = {5'd26, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 25 {'a': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 25, 'op': 'read'}
    instructions[3320] = {5'd0, 4'd2, 4'd0, 16'd540};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 25 {'literal': 540, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 25, 'op': 'literal'}
    instructions[3321] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 25 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 25, 'op': 'store'}
    instructions[3322] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 25 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 25, 'op': 'addl'}
    instructions[3323] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 25 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 25, 'op': 'addl'}
    instructions[3324] = {5'd16, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 25 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 25, 'op': 'return'}
    instructions[3325] = {5'd1, 4'd3, 4'd3, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 78 {'a': 3, 'literal': 3, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 78, 'op': 'addl'}
    instructions[3326] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 84 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 84, 'op': 'literal'}
    instructions[3327] = {5'd1, 4'd2, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 84 {'a': 4, 'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 84, 'op': 'addl'}
    instructions[3328] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 84 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 84, 'op': 'store'}
    instructions[3329] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 85 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 85, 'op': 'addl'}
    instructions[3330] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 85 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 85, 'op': 'addl'}
    instructions[3331] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 85 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 85, 'op': 'load'}
    instructions[3332] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 85 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 85, 'op': 'store'}
    instructions[3333] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 85 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 85, 'op': 'addl'}
    instructions[3334] = {5'd1, 4'd8, 4'd4, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 85 {'a': 4, 'literal': -2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 85, 'op': 'addl'}
    instructions[3335] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 85 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 85, 'op': 'addl'}
    instructions[3336] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 85 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 85, 'op': 'load'}
    instructions[3337] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 85 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 85, 'op': 'store'}
    instructions[3338] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 85 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 85, 'op': 'addl'}
    instructions[3339] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 85 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 85, 'op': 'literal'}
    instructions[3340] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 85 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 85, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3341] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 85 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 85, 'op': 'load'}
    instructions[3342] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 85 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 85, 'op': 'add'}
    instructions[3343] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 85 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 85, 'op': 'addl'}
    instructions[3344] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 85 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 85, 'op': 'load'}
    instructions[3345] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 85 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 85, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3346] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 85 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 85, 'op': 'load'}
    instructions[3347] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 85 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 85, 'op': 'add'}
    instructions[3348] = {5'd1, 4'd2, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 85 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 85, 'op': 'addl'}
    instructions[3349] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 85 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 85, 'op': 'store'}
    instructions[3350] = {5'd1, 4'd8, 4'd4, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 86 {'a': 4, 'literal': -2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 86, 'op': 'addl'}
    instructions[3351] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 86 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 86, 'op': 'addl'}
    instructions[3352] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 86 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 86, 'op': 'load'}
    instructions[3353] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 86 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 86, 'op': 'store'}
    instructions[3354] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 86 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 86, 'op': 'addl'}
    instructions[3355] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 86 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 86, 'op': 'literal'}
    instructions[3356] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 86 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 86, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3357] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 86 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 86, 'op': 'load'}
    instructions[3358] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 86 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 86, 'op': 'add'}
    instructions[3359] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 86 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 86, 'op': 'addl'}
    instructions[3360] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 86 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 86, 'op': 'load'}
    instructions[3361] = {5'd1, 4'd2, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 86 {'a': 4, 'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 86, 'op': 'addl'}
    instructions[3362] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 86 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 86, 'op': 'store'}
    instructions[3363] = {5'd0, 4'd8, 4'd0, 16'd65535};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 87 {'literal': 65535, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 87, 'op': 'literal'}
    instructions[3364] = {5'd3, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 87 {'a': 8, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 87, 'op': 'literal_hi'}
    instructions[3365] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 87 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 87, 'op': 'store'}
    instructions[3366] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 87 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 87, 'op': 'addl'}
    instructions[3367] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 87 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 87, 'op': 'addl'}
    instructions[3368] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 87 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 87, 'op': 'addl'}
    instructions[3369] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 87 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 87, 'op': 'load'}
    instructions[3370] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 87 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 87, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3371] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 87 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 87, 'op': 'load'}
    instructions[3372] = {5'd19, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 87 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 87, 'op': 'unsigned_greater'}
    instructions[3373] = {5'd8, 4'd0, 4'd8, 16'd3386};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 87 {'a': 8, 'label': 3386, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 87, 'op': 'jmp_if_false'}
    instructions[3374] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 87 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 87, 'op': 'literal'}
    instructions[3375] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 87 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 87, 'op': 'store'}
    instructions[3376] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 87 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 87, 'op': 'addl'}
    instructions[3377] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 87 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 87, 'op': 'addl'}
    instructions[3378] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 87 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 87, 'op': 'addl'}
    instructions[3379] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 87 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 87, 'op': 'load'}
    instructions[3380] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 87 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 87, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3381] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 87 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 87, 'op': 'load'}
    instructions[3382] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 87 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 87, 'op': 'add'}
    instructions[3383] = {5'd1, 4'd2, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 87 {'a': 4, 'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 87, 'op': 'addl'}
    instructions[3384] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 87 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 87, 'op': 'store'}
    instructions[3385] = {5'd10, 4'd0, 4'd0, 16'd3386};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 87 {'label': 3386, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 87, 'op': 'goto'}
    instructions[3386] = {5'd1, 4'd8, 4'd4, -16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90 {'a': 4, 'literal': -3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90, 'op': 'addl'}
    instructions[3387] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90, 'op': 'addl'}
    instructions[3388] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90, 'op': 'load'}
    instructions[3389] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90, 'op': 'store'}
    instructions[3390] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90, 'op': 'addl'}
    instructions[3391] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90, 'op': 'literal'}
    instructions[3392] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3393] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90, 'op': 'load'}
    instructions[3394] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90, 'op': 'add'}
    instructions[3395] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90, 'op': 'addl'}
    instructions[3396] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90, 'op': 'load'}
    instructions[3397] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90, 'op': 'store'}
    instructions[3398] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90, 'op': 'addl'}
    instructions[3399] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90, 'op': 'addl'}
    instructions[3400] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90, 'op': 'addl'}
    instructions[3401] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90, 'op': 'load'}
    instructions[3402] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3403] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90, 'op': 'load'}
    instructions[3404] = {5'd13, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90, 'op': 'not_equal'}
    instructions[3405] = {5'd12, 4'd0, 4'd8, 16'd3425};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90 {'a': 8, 'label': 3425, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90, 'op': 'jmp_if_true'}
    instructions[3406] = {5'd1, 4'd8, 4'd4, -16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90 {'a': 4, 'literal': -3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90, 'op': 'addl'}
    instructions[3407] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90, 'op': 'addl'}
    instructions[3408] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90, 'op': 'load'}
    instructions[3409] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90, 'op': 'store'}
    instructions[3410] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90, 'op': 'addl'}
    instructions[3411] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90, 'op': 'literal'}
    instructions[3412] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3413] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90, 'op': 'load'}
    instructions[3414] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90, 'op': 'add'}
    instructions[3415] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90, 'op': 'addl'}
    instructions[3416] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90, 'op': 'load'}
    instructions[3417] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90, 'op': 'store'}
    instructions[3418] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90, 'op': 'addl'}
    instructions[3419] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90, 'op': 'addl'}
    instructions[3420] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90, 'op': 'addl'}
    instructions[3421] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90, 'op': 'load'}
    instructions[3422] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3423] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90, 'op': 'load'}
    instructions[3424] = {5'd13, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90, 'op': 'not_equal'}
    instructions[3425] = {5'd8, 4'd0, 4'd8, 16'd3466};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90 {'a': 8, 'label': 3466, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90, 'op': 'jmp_if_false'}
    instructions[3426] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 91 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 91, 'op': 'addl'}
    instructions[3427] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 91 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 91, 'op': 'addl'}
    instructions[3428] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 91 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 91, 'op': 'load'}
    instructions[3429] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 91 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 91, 'op': 'store'}
    instructions[3430] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 91 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 91, 'op': 'addl'}
    instructions[3431] = {5'd1, 4'd8, 4'd4, -16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 91 {'a': 4, 'literal': -3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 91, 'op': 'addl'}
    instructions[3432] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 91 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 91, 'op': 'addl'}
    instructions[3433] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 91 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 91, 'op': 'load'}
    instructions[3434] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 91 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 91, 'op': 'store'}
    instructions[3435] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 91 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 91, 'op': 'addl'}
    instructions[3436] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 91 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 91, 'op': 'literal'}
    instructions[3437] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 91 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 91, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3438] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 91 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 91, 'op': 'load'}
    instructions[3439] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 91 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 91, 'op': 'add'}
    instructions[3440] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 91 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 91, 'op': 'addl'}
    instructions[3441] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 91 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 91, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3442] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 91 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 91, 'op': 'load'}
    instructions[3443] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 91 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 91, 'op': 'store'}
    instructions[3444] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 92 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 92, 'op': 'addl'}
    instructions[3445] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 92 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 92, 'op': 'addl'}
    instructions[3446] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 92 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 92, 'op': 'load'}
    instructions[3447] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 92 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 92, 'op': 'store'}
    instructions[3448] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 92 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 92, 'op': 'addl'}
    instructions[3449] = {5'd1, 4'd8, 4'd4, -16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 92 {'a': 4, 'literal': -3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 92, 'op': 'addl'}
    instructions[3450] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 92 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 92, 'op': 'addl'}
    instructions[3451] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 92 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 92, 'op': 'load'}
    instructions[3452] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 92 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 92, 'op': 'store'}
    instructions[3453] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 92 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 92, 'op': 'addl'}
    instructions[3454] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 92 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 92, 'op': 'literal'}
    instructions[3455] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 92 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 92, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3456] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 92 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 92, 'op': 'load'}
    instructions[3457] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 92 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 92, 'op': 'add'}
    instructions[3458] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 92 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 92, 'op': 'addl'}
    instructions[3459] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 92 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 92, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3460] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 92 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 92, 'op': 'load'}
    instructions[3461] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 92 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 92, 'op': 'store'}
    instructions[3462] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 93 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 93, 'op': 'literal'}
    instructions[3463] = {5'd1, 4'd2, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 93 {'a': 4, 'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 93, 'op': 'addl'}
    instructions[3464] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 93 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 93, 'op': 'store'}
    instructions[3465] = {5'd10, 4'd0, 4'd0, 16'd3466};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90 {'label': 3466, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 90, 'op': 'goto'}
    instructions[3466] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 95 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 95, 'op': 'addl'}
    instructions[3467] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 95 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 95, 'op': 'addl'}
    instructions[3468] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 95 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 95, 'op': 'load'}
    instructions[3469] = {5'd0, 4'd2, 4'd0, 16'd582};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 95 {'literal': 582, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 95, 'op': 'literal'}
    instructions[3470] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 95 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 95, 'op': 'store'}
    instructions[3471] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 95 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 95, 'op': 'addl'}
    instructions[3472] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 95 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 95, 'op': 'addl'}
    instructions[3473] = {5'd16, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 95 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 95, 'op': 'return'}
    instructions[3474] = {5'd1, 4'd3, 4'd3, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 492 {'a': 3, 'literal': 3, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 492, 'op': 'addl'}
    instructions[3475] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 495 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 495, 'op': 'literal'}
    instructions[3476] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 495 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 495, 'op': 'store'}
    instructions[3477] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 495 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 495, 'op': 'addl'}
    instructions[3478] = {5'd0, 4'd8, 4'd0, 16'd16};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 495 {'literal': 16, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 495, 'op': 'literal'}
    instructions[3479] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 495 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 495, 'op': 'addl'}
    instructions[3480] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 495 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 495, 'op': 'load'}
    instructions[3481] = {5'd14, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 495 {'a': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 495, 'op': 'ready'}
    instructions[3482] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 495 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 495, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3483] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 495 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 495, 'op': 'load'}
    instructions[3484] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 495 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 495, 'op': 'equal'}
    instructions[3485] = {5'd8, 4'd0, 4'd8, 16'd3493};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 495 {'a': 8, 'label': 3493, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 495, 'op': 'jmp_if_false'}
    instructions[3486] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 496 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 496, 'op': 'literal'}
    instructions[3487] = {5'd0, 4'd2, 4'd0, 16'd543};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 496 {'literal': 543, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 496, 'op': 'literal'}
    instructions[3488] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 496 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 496, 'op': 'store'}
    instructions[3489] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 496 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 496, 'op': 'addl'}
    instructions[3490] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 496 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 496, 'op': 'addl'}
    instructions[3491] = {5'd16, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 496 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 496, 'op': 'return'}
    instructions[3492] = {5'd10, 4'd0, 4'd0, 16'd3493};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 495 {'label': 3493, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 495, 'op': 'goto'}
    instructions[3493] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 499 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 499, 'op': 'addl'}
    instructions[3494] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 499 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 499, 'op': 'addl'}
    instructions[3495] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 499 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 499, 'op': 'load'}
    instructions[3496] = {5'd1, 4'd2, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 499 {'a': 4, 'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 499, 'op': 'addl'}
    instructions[3497] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 499 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 499, 'op': 'store'}
    instructions[3498] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 500 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 500, 'op': 'store'}
    instructions[3499] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 500 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 500, 'op': 'addl'}
    instructions[3500] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 500 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 500, 'op': 'store'}
    instructions[3501] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 500 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 500, 'op': 'addl'}
    instructions[3502] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 500 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 500, 'op': 'addl'}
    instructions[3503] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 500 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 500, 'op': 'addl'}
    instructions[3504] = {5'd4, 4'd6, 4'd0, 16'd3598};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 500 {'z': 6, 'label': 3598, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 500, 'op': 'call'}
    instructions[3505] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 500 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 500, 'op': 'addl'}
    instructions[3506] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 500 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 500, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3507] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 500 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 500, 'op': 'load'}
    instructions[3508] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 500 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 500, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3509] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 500 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 500, 'op': 'load'}
    instructions[3510] = {5'd0, 4'd2, 4'd0, 16'd584};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 500 {'literal': 584, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 500, 'op': 'literal'}
    instructions[3511] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 500 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 500, 'op': 'load'}
    instructions[3512] = {5'd1, 4'd2, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 500 {'a': 4, 'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 500, 'op': 'addl'}
    instructions[3513] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 500 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 500, 'op': 'store'}
    instructions[3514] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501, 'op': 'literal'}
    instructions[3515] = {5'd1, 4'd2, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501, 'op': 'addl'}
    instructions[3516] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501, 'op': 'store'}
    instructions[3517] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501, 'op': 'addl'}
    instructions[3518] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501, 'op': 'addl'}
    instructions[3519] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501, 'op': 'load'}
    instructions[3520] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501, 'op': 'store'}
    instructions[3521] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501, 'op': 'addl'}
    instructions[3522] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501, 'op': 'addl'}
    instructions[3523] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501, 'op': 'addl'}
    instructions[3524] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501, 'op': 'load'}
    instructions[3525] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3526] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501, 'op': 'load'}
    instructions[3527] = {5'd19, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501, 'op': 'unsigned_greater'}
    instructions[3528] = {5'd8, 4'd0, 4'd8, 16'd3590};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501 {'a': 8, 'label': 3590, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501, 'op': 'jmp_if_false'}
    instructions[3529] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502, 'op': 'store'}
    instructions[3530] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502, 'op': 'addl'}
    instructions[3531] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502, 'op': 'store'}
    instructions[3532] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502, 'op': 'addl'}
    instructions[3533] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502, 'op': 'addl'}
    instructions[3534] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502, 'op': 'addl'}
    instructions[3535] = {5'd4, 4'd6, 4'd0, 16'd3598};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502 {'z': 6, 'label': 3598, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502, 'op': 'call'}
    instructions[3536] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502, 'op': 'addl'}
    instructions[3537] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3538] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502, 'op': 'load'}
    instructions[3539] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3540] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502, 'op': 'load'}
    instructions[3541] = {5'd0, 4'd2, 4'd0, 16'd584};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502 {'literal': 584, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502, 'op': 'literal'}
    instructions[3542] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502, 'op': 'load'}
    instructions[3543] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502, 'op': 'store'}
    instructions[3544] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502, 'op': 'addl'}
    instructions[3545] = {5'd1, 4'd8, 4'd4, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502 {'a': 4, 'literal': -2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502, 'op': 'addl'}
    instructions[3546] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502, 'op': 'addl'}
    instructions[3547] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502, 'op': 'load'}
    instructions[3548] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502, 'op': 'store'}
    instructions[3549] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502, 'op': 'addl'}
    instructions[3550] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502, 'op': 'addl'}
    instructions[3551] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502, 'op': 'addl'}
    instructions[3552] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502, 'op': 'load'}
    instructions[3553] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3554] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502, 'op': 'load'}
    instructions[3555] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502, 'op': 'add'}
    instructions[3556] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502, 'op': 'addl'}
    instructions[3557] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3558] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502, 'op': 'load'}
    instructions[3559] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 502, 'op': 'store'}
    instructions[3560] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 503 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 503, 'op': 'addl'}
    instructions[3561] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 503 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 503, 'op': 'addl'}
    instructions[3562] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 503 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 503, 'op': 'load'}
    instructions[3563] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 503 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 503, 'op': 'store'}
    instructions[3564] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 503 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 503, 'op': 'addl'}
    instructions[3565] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 503 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 503, 'op': 'literal'}
    instructions[3566] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 503 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 503, 'op': 'store'}
    instructions[3567] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 503 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 503, 'op': 'addl'}
    instructions[3568] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 503 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 503, 'op': 'addl'}
    instructions[3569] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 503 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 503, 'op': 'addl'}
    instructions[3570] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 503 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 503, 'op': 'load'}
    instructions[3571] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 503 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 503, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3572] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 503 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 503, 'op': 'load'}
    instructions[3573] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 503 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 503, 'op': 'add'}
    instructions[3574] = {5'd1, 4'd2, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 503 {'a': 4, 'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 503, 'op': 'addl'}
    instructions[3575] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 503 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 503, 'op': 'store'}
    instructions[3576] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 503 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 503, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3577] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 503 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 503, 'op': 'load'}
    instructions[3578] = {5'd0, 4'd8, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501 {'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501, 'op': 'literal'}
    instructions[3579] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501, 'op': 'store'}
    instructions[3580] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501, 'op': 'addl'}
    instructions[3581] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501, 'op': 'addl'}
    instructions[3582] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501, 'op': 'addl'}
    instructions[3583] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501, 'op': 'load'}
    instructions[3584] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3585] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501, 'op': 'load'}
    instructions[3586] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501, 'op': 'add'}
    instructions[3587] = {5'd1, 4'd2, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501, 'op': 'addl'}
    instructions[3588] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501, 'op': 'store'}
    instructions[3589] = {5'd10, 4'd0, 4'd0, 16'd3517};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501 {'label': 3517, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 501, 'op': 'goto'}
    instructions[3590] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 505 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 505, 'op': 'addl'}
    instructions[3591] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 505 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 505, 'op': 'addl'}
    instructions[3592] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 505 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 505, 'op': 'load'}
    instructions[3593] = {5'd0, 4'd2, 4'd0, 16'd543};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 505 {'literal': 543, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 505, 'op': 'literal'}
    instructions[3594] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 505 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 505, 'op': 'store'}
    instructions[3595] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 505 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 505, 'op': 'addl'}
    instructions[3596] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 505 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 505, 'op': 'addl'}
    instructions[3597] = {5'd16, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 505 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 505, 'op': 'return'}
    instructions[3598] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 30 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 30, 'op': 'addl'}
    instructions[3599] = {5'd0, 4'd8, 4'd0, 16'd16};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 31 {'literal': 16, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 31, 'op': 'literal'}
    instructions[3600] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 31 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 31, 'op': 'addl'}
    instructions[3601] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 31 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 31, 'op': 'load'}
    instructions[3602] = {5'd26, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 31 {'a': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 31, 'op': 'read'}
    instructions[3603] = {5'd0, 4'd2, 4'd0, 16'd584};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 31 {'literal': 584, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 31, 'op': 'literal'}
    instructions[3604] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 31 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 31, 'op': 'store'}
    instructions[3605] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 31 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 31, 'op': 'addl'}
    instructions[3606] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 31 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 31, 'op': 'addl'}
    instructions[3607] = {5'd16, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 31 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 31, 'op': 'return'}
    instructions[3608] = {5'd1, 4'd3, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 445 {'a': 3, 'literal': 7, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 445, 'op': 'addl'}
    instructions[3609] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 449 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 449, 'op': 'store'}
    instructions[3610] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 449 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 449, 'op': 'addl'}
    instructions[3611] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 449 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 449, 'op': 'store'}
    instructions[3612] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 449 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 449, 'op': 'addl'}
    instructions[3613] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 449 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 449, 'op': 'addl'}
    instructions[3614] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 449 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 449, 'op': 'addl'}
    instructions[3615] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 449 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 449, 'op': 'load'}
    instructions[3616] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 449 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 449, 'op': 'store'}
    instructions[3617] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 449 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 449, 'op': 'addl'}
    instructions[3618] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 449 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 449, 'op': 'addl'}
    instructions[3619] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 449 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 449, 'op': 'addl'}
    instructions[3620] = {5'd4, 4'd6, 4'd0, 16'd4131};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 449 {'z': 6, 'label': 4131, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 449, 'op': 'call'}
    instructions[3621] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 449 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 449, 'op': 'addl'}
    instructions[3622] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 449 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 449, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3623] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 449 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 449, 'op': 'load'}
    instructions[3624] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 449 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 449, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3625] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 449 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 449, 'op': 'load'}
    instructions[3626] = {5'd0, 4'd2, 4'd0, 16'd17};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 449 {'literal': 17, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 449, 'op': 'literal'}
    instructions[3627] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 449 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 449, 'op': 'load'}
    instructions[3628] = {5'd1, 4'd2, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 449 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 449, 'op': 'addl'}
    instructions[3629] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 449 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 449, 'op': 'store'}
    instructions[3630] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452, 'op': 'literal'}
    instructions[3631] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452, 'op': 'store'}
    instructions[3632] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452, 'op': 'addl'}
    instructions[3633] = {5'd0, 4'd8, 4'd0, 16'd15};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452 {'literal': 15, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452, 'op': 'literal'}
    instructions[3634] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452, 'op': 'store'}
    instructions[3635] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452, 'op': 'addl'}
    instructions[3636] = {5'd0, 4'd8, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452 {'literal': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452, 'op': 'literal'}
    instructions[3637] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452, 'op': 'store'}
    instructions[3638] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452, 'op': 'addl'}
    instructions[3639] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452, 'op': 'addl'}
    instructions[3640] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452, 'op': 'addl'}
    instructions[3641] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452, 'op': 'load'}
    instructions[3642] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452, 'op': 'store'}
    instructions[3643] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452, 'op': 'addl'}
    instructions[3644] = {5'd0, 4'd8, 4'd0, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452 {'literal': 7, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452, 'op': 'literal'}
    instructions[3645] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3646] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452, 'op': 'load'}
    instructions[3647] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452, 'op': 'add'}
    instructions[3648] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452, 'op': 'addl'}
    instructions[3649] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452, 'op': 'load'}
    instructions[3650] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3651] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452, 'op': 'load'}
    instructions[3652] = {5'd27, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452, 'op': 'shift_right'}
    instructions[3653] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3654] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452, 'op': 'load'}
    instructions[3655] = {5'd22, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452, 'op': 'and'}
    instructions[3656] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3657] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452, 'op': 'load'}
    instructions[3658] = {5'd28, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452, 'op': 'shift_left'}
    instructions[3659] = {5'd1, 4'd2, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452 {'a': 4, 'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452, 'op': 'addl'}
    instructions[3660] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 452, 'op': 'store'}
    instructions[3661] = {5'd0, 4'd8, 4'd0, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 453 {'literal': 7, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 453, 'op': 'literal'}
    instructions[3662] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 453 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 453, 'op': 'store'}
    instructions[3663] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 453 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 453, 'op': 'addl'}
    instructions[3664] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 453 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 453, 'op': 'addl'}
    instructions[3665] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 453 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 453, 'op': 'addl'}
    instructions[3666] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 453 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 453, 'op': 'load'}
    instructions[3667] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 453 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 453, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3668] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 453 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 453, 'op': 'load'}
    instructions[3669] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 453 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 453, 'op': 'add'}
    instructions[3670] = {5'd1, 4'd2, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 453 {'a': 4, 'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 453, 'op': 'addl'}
    instructions[3671] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 453 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 453, 'op': 'store'}
    instructions[3672] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 455 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 455, 'op': 'addl'}
    instructions[3673] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 455 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 455, 'op': 'addl'}
    instructions[3674] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 455 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 455, 'op': 'load'}
    instructions[3675] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 455 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 455, 'op': 'store'}
    instructions[3676] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 455 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 455, 'op': 'addl'}
    instructions[3677] = {5'd0, 4'd8, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 455 {'literal': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 455, 'op': 'literal'}
    instructions[3678] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 455 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 455, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3679] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 455 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 455, 'op': 'load'}
    instructions[3680] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 455 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 455, 'op': 'add'}
    instructions[3681] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 455 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 455, 'op': 'addl'}
    instructions[3682] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 455 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 455, 'op': 'load'}
    instructions[3683] = {5'd1, 4'd2, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 455 {'a': 4, 'literal': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 455, 'op': 'addl'}
    instructions[3684] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 455 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 455, 'op': 'store'}
    instructions[3685] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 456 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 456, 'op': 'literal'}
    instructions[3686] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 456 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 456, 'op': 'store'}
    instructions[3687] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 456 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 456, 'op': 'addl'}
    instructions[3688] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 456 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 456, 'op': 'addl'}
    instructions[3689] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 456 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 456, 'op': 'addl'}
    instructions[3690] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 456 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 456, 'op': 'load'}
    instructions[3691] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 456 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 456, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3692] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 456 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 456, 'op': 'load'}
    instructions[3693] = {5'd28, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 456 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 456, 'op': 'shift_left'}
    instructions[3694] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 456 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 456, 'op': 'store'}
    instructions[3695] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 456 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 456, 'op': 'addl'}
    instructions[3696] = {5'd1, 4'd8, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 456 {'a': 4, 'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 456, 'op': 'addl'}
    instructions[3697] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 456 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 456, 'op': 'addl'}
    instructions[3698] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 456 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 456, 'op': 'load'}
    instructions[3699] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 456 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 456, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3700] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 456 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 456, 'op': 'load'}
    instructions[3701] = {5'd9, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 456 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 456, 'op': 'subtract'}
    instructions[3702] = {5'd1, 4'd2, 4'd4, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 456 {'a': 4, 'literal': 4, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 456, 'op': 'addl'}
    instructions[3703] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 456 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 456, 'op': 'store'}
    instructions[3704] = {5'd0, 4'd8, 4'd0, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457 {'literal': 10, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457, 'op': 'literal'}
    instructions[3705] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457, 'op': 'store'}
    instructions[3706] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457, 'op': 'addl'}
    instructions[3707] = {5'd0, 4'd8, 4'd0, 16'd61440};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457 {'literal': 61440, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457, 'op': 'literal'}
    instructions[3708] = {5'd3, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457 {'a': 8, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457, 'op': 'literal_hi'}
    instructions[3709] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457, 'op': 'store'}
    instructions[3710] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457, 'op': 'addl'}
    instructions[3711] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457, 'op': 'addl'}
    instructions[3712] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457, 'op': 'addl'}
    instructions[3713] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457, 'op': 'load'}
    instructions[3714] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457, 'op': 'store'}
    instructions[3715] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457, 'op': 'addl'}
    instructions[3716] = {5'd0, 4'd8, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457 {'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457, 'op': 'literal'}
    instructions[3717] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457, 'op': 'store'}
    instructions[3718] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457, 'op': 'addl'}
    instructions[3719] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457, 'op': 'addl'}
    instructions[3720] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457, 'op': 'addl'}
    instructions[3721] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457, 'op': 'load'}
    instructions[3722] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3723] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457, 'op': 'load'}
    instructions[3724] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457, 'op': 'add'}
    instructions[3725] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3726] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457, 'op': 'load'}
    instructions[3727] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457, 'op': 'add'}
    instructions[3728] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457, 'op': 'addl'}
    instructions[3729] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457, 'op': 'load'}
    instructions[3730] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3731] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457, 'op': 'load'}
    instructions[3732] = {5'd22, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457, 'op': 'and'}
    instructions[3733] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3734] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457, 'op': 'load'}
    instructions[3735] = {5'd18, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457, 'op': 'unsigned_shift_right'}
    instructions[3736] = {5'd1, 4'd2, 4'd4, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457 {'a': 4, 'literal': 6, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457, 'op': 'addl'}
    instructions[3737] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 457, 'op': 'store'}
    instructions[3738] = {5'd1, 4'd8, 4'd4, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 458 {'a': 4, 'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 458, 'op': 'addl'}
    instructions[3739] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 458 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 458, 'op': 'addl'}
    instructions[3740] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 458 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 458, 'op': 'load'}
    instructions[3741] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 458 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 458, 'op': 'store'}
    instructions[3742] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 458 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 458, 'op': 'addl'}
    instructions[3743] = {5'd1, 4'd8, 4'd4, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 458 {'a': 4, 'literal': 4, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 458, 'op': 'addl'}
    instructions[3744] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 458 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 458, 'op': 'addl'}
    instructions[3745] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 458 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 458, 'op': 'load'}
    instructions[3746] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 458 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 458, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3747] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 458 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 458, 'op': 'load'}
    instructions[3748] = {5'd9, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 458 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 458, 'op': 'subtract'}
    instructions[3749] = {5'd0, 4'd2, 4'd0, 16'd581};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 458 {'literal': 581, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 458, 'op': 'literal'}
    instructions[3750] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 458 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 458, 'op': 'store'}
    instructions[3751] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 459 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 459, 'op': 'literal'}
    instructions[3752] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 459 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 459, 'op': 'store'}
    instructions[3753] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 459 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 459, 'op': 'addl'}
    instructions[3754] = {5'd1, 4'd8, 4'd4, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 459 {'a': 4, 'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 459, 'op': 'addl'}
    instructions[3755] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 459 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 459, 'op': 'addl'}
    instructions[3756] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 459 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 459, 'op': 'load'}
    instructions[3757] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 459 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 459, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3758] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 459 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 459, 'op': 'load'}
    instructions[3759] = {5'd18, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 459 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 459, 'op': 'unsigned_shift_right'}
    instructions[3760] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 459 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 459, 'op': 'store'}
    instructions[3761] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 459 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 459, 'op': 'addl'}
    instructions[3762] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 459 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 459, 'op': 'addl'}
    instructions[3763] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 459 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 459, 'op': 'addl'}
    instructions[3764] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 459 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 459, 'op': 'load'}
    instructions[3765] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 459 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 459, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3766] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 459 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 459, 'op': 'load'}
    instructions[3767] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 459 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 459, 'op': 'add'}
    instructions[3768] = {5'd0, 4'd2, 4'd0, 16'd21};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 459 {'literal': 21, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 459, 'op': 'literal'}
    instructions[3769] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 459 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 459, 'op': 'store'}
    instructions[3770] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 462 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 462, 'op': 'addl'}
    instructions[3771] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 462 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 462, 'op': 'addl'}
    instructions[3772] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 462 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 462, 'op': 'load'}
    instructions[3773] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 462 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 462, 'op': 'store'}
    instructions[3774] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 462 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 462, 'op': 'addl'}
    instructions[3775] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 462 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 462, 'op': 'literal'}
    instructions[3776] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 462 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 462, 'op': 'store'}
    instructions[3777] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 462 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 462, 'op': 'addl'}
    instructions[3778] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 462 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 462, 'op': 'addl'}
    instructions[3779] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 462 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 462, 'op': 'addl'}
    instructions[3780] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 462 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 462, 'op': 'load'}
    instructions[3781] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 462 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 462, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3782] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 462 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 462, 'op': 'load'}
    instructions[3783] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 462 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 462, 'op': 'add'}
    instructions[3784] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 462 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 462, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3785] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 462 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 462, 'op': 'load'}
    instructions[3786] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 462 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 462, 'op': 'add'}
    instructions[3787] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 462 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 462, 'op': 'addl'}
    instructions[3788] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 462 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 462, 'op': 'load'}
    instructions[3789] = {5'd0, 4'd2, 4'd0, 16'd651};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 462 {'literal': 651, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 462, 'op': 'literal'}
    instructions[3790] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 462 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 462, 'op': 'store'}
    instructions[3791] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 463 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 463, 'op': 'addl'}
    instructions[3792] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 463 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 463, 'op': 'addl'}
    instructions[3793] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 463 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 463, 'op': 'load'}
    instructions[3794] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 463 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 463, 'op': 'store'}
    instructions[3795] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 463 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 463, 'op': 'addl'}
    instructions[3796] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 463 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 463, 'op': 'literal'}
    instructions[3797] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 463 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 463, 'op': 'store'}
    instructions[3798] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 463 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 463, 'op': 'addl'}
    instructions[3799] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 463 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 463, 'op': 'addl'}
    instructions[3800] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 463 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 463, 'op': 'addl'}
    instructions[3801] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 463 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 463, 'op': 'load'}
    instructions[3802] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 463 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 463, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3803] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 463 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 463, 'op': 'load'}
    instructions[3804] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 463 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 463, 'op': 'add'}
    instructions[3805] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 463 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 463, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3806] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 463 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 463, 'op': 'load'}
    instructions[3807] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 463 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 463, 'op': 'add'}
    instructions[3808] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 463 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 463, 'op': 'addl'}
    instructions[3809] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 463 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 463, 'op': 'load'}
    instructions[3810] = {5'd0, 4'd2, 4'd0, 16'd628};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 463 {'literal': 628, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 463, 'op': 'literal'}
    instructions[3811] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 463 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 463, 'op': 'store'}
    instructions[3812] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464, 'op': 'addl'}
    instructions[3813] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464, 'op': 'addl'}
    instructions[3814] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464, 'op': 'load'}
    instructions[3815] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464, 'op': 'store'}
    instructions[3816] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464, 'op': 'addl'}
    instructions[3817] = {5'd0, 4'd8, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464 {'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464, 'op': 'literal'}
    instructions[3818] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464, 'op': 'store'}
    instructions[3819] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464, 'op': 'addl'}
    instructions[3820] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464, 'op': 'addl'}
    instructions[3821] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464, 'op': 'addl'}
    instructions[3822] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464, 'op': 'load'}
    instructions[3823] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3824] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464, 'op': 'load'}
    instructions[3825] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464, 'op': 'add'}
    instructions[3826] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3827] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464, 'op': 'load'}
    instructions[3828] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464, 'op': 'add'}
    instructions[3829] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464, 'op': 'addl'}
    instructions[3830] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464, 'op': 'load'}
    instructions[3831] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464, 'op': 'store'}
    instructions[3832] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464, 'op': 'addl'}
    instructions[3833] = {5'd0, 4'd8, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464 {'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464, 'op': 'literal'}
    instructions[3834] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464, 'op': 'store'}
    instructions[3835] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464, 'op': 'addl'}
    instructions[3836] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464, 'op': 'literal'}
    instructions[3837] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3838] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464, 'op': 'load'}
    instructions[3839] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464, 'op': 'add'}
    instructions[3840] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464, 'op': 'addl'}
    instructions[3841] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3842] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464, 'op': 'load'}
    instructions[3843] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 464, 'op': 'store'}
    instructions[3844] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465, 'op': 'addl'}
    instructions[3845] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465, 'op': 'addl'}
    instructions[3846] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465, 'op': 'load'}
    instructions[3847] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465, 'op': 'store'}
    instructions[3848] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465, 'op': 'addl'}
    instructions[3849] = {5'd0, 4'd8, 4'd0, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465 {'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465, 'op': 'literal'}
    instructions[3850] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465, 'op': 'store'}
    instructions[3851] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465, 'op': 'addl'}
    instructions[3852] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465, 'op': 'addl'}
    instructions[3853] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465, 'op': 'addl'}
    instructions[3854] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465, 'op': 'load'}
    instructions[3855] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3856] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465, 'op': 'load'}
    instructions[3857] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465, 'op': 'add'}
    instructions[3858] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3859] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465, 'op': 'load'}
    instructions[3860] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465, 'op': 'add'}
    instructions[3861] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465, 'op': 'addl'}
    instructions[3862] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465, 'op': 'load'}
    instructions[3863] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465, 'op': 'store'}
    instructions[3864] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465, 'op': 'addl'}
    instructions[3865] = {5'd0, 4'd8, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465 {'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465, 'op': 'literal'}
    instructions[3866] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465, 'op': 'store'}
    instructions[3867] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465, 'op': 'addl'}
    instructions[3868] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465, 'op': 'literal'}
    instructions[3869] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3870] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465, 'op': 'load'}
    instructions[3871] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465, 'op': 'add'}
    instructions[3872] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465, 'op': 'addl'}
    instructions[3873] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3874] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465, 'op': 'load'}
    instructions[3875] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 465, 'op': 'store'}
    instructions[3876] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466, 'op': 'addl'}
    instructions[3877] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466, 'op': 'addl'}
    instructions[3878] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466, 'op': 'load'}
    instructions[3879] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466, 'op': 'store'}
    instructions[3880] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466, 'op': 'addl'}
    instructions[3881] = {5'd0, 4'd8, 4'd0, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466 {'literal': 4, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466, 'op': 'literal'}
    instructions[3882] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466, 'op': 'store'}
    instructions[3883] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466, 'op': 'addl'}
    instructions[3884] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466, 'op': 'addl'}
    instructions[3885] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466, 'op': 'addl'}
    instructions[3886] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466, 'op': 'load'}
    instructions[3887] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3888] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466, 'op': 'load'}
    instructions[3889] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466, 'op': 'add'}
    instructions[3890] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3891] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466, 'op': 'load'}
    instructions[3892] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466, 'op': 'add'}
    instructions[3893] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466, 'op': 'addl'}
    instructions[3894] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466, 'op': 'load'}
    instructions[3895] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466, 'op': 'store'}
    instructions[3896] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466, 'op': 'addl'}
    instructions[3897] = {5'd0, 4'd8, 4'd0, 16'd18};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466 {'literal': 18, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466, 'op': 'literal'}
    instructions[3898] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466, 'op': 'store'}
    instructions[3899] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466, 'op': 'addl'}
    instructions[3900] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466, 'op': 'literal'}
    instructions[3901] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3902] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466, 'op': 'load'}
    instructions[3903] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466, 'op': 'add'}
    instructions[3904] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466, 'op': 'addl'}
    instructions[3905] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3906] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466, 'op': 'load'}
    instructions[3907] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 466, 'op': 'store'}
    instructions[3908] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467, 'op': 'addl'}
    instructions[3909] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467, 'op': 'addl'}
    instructions[3910] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467, 'op': 'load'}
    instructions[3911] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467, 'op': 'store'}
    instructions[3912] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467, 'op': 'addl'}
    instructions[3913] = {5'd0, 4'd8, 4'd0, 16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467 {'literal': 5, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467, 'op': 'literal'}
    instructions[3914] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467, 'op': 'store'}
    instructions[3915] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467, 'op': 'addl'}
    instructions[3916] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467, 'op': 'addl'}
    instructions[3917] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467, 'op': 'addl'}
    instructions[3918] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467, 'op': 'load'}
    instructions[3919] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3920] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467, 'op': 'load'}
    instructions[3921] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467, 'op': 'add'}
    instructions[3922] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3923] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467, 'op': 'load'}
    instructions[3924] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467, 'op': 'add'}
    instructions[3925] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467, 'op': 'addl'}
    instructions[3926] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467, 'op': 'load'}
    instructions[3927] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467, 'op': 'store'}
    instructions[3928] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467, 'op': 'addl'}
    instructions[3929] = {5'd0, 4'd8, 4'd0, 16'd18};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467 {'literal': 18, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467, 'op': 'literal'}
    instructions[3930] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467, 'op': 'store'}
    instructions[3931] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467, 'op': 'addl'}
    instructions[3932] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467, 'op': 'literal'}
    instructions[3933] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3934] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467, 'op': 'load'}
    instructions[3935] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467, 'op': 'add'}
    instructions[3936] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467, 'op': 'addl'}
    instructions[3937] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3938] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467, 'op': 'load'}
    instructions[3939] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 467, 'op': 'store'}
    instructions[3940] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 468 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 468, 'op': 'addl'}
    instructions[3941] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 468 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 468, 'op': 'addl'}
    instructions[3942] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 468 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 468, 'op': 'load'}
    instructions[3943] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 468 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 468, 'op': 'store'}
    instructions[3944] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 468 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 468, 'op': 'addl'}
    instructions[3945] = {5'd0, 4'd8, 4'd0, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 468 {'literal': 7, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 468, 'op': 'literal'}
    instructions[3946] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 468 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 468, 'op': 'store'}
    instructions[3947] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 468 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 468, 'op': 'addl'}
    instructions[3948] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 468 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 468, 'op': 'addl'}
    instructions[3949] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 468 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 468, 'op': 'addl'}
    instructions[3950] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 468 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 468, 'op': 'load'}
    instructions[3951] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 468 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 468, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3952] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 468 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 468, 'op': 'load'}
    instructions[3953] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 468 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 468, 'op': 'add'}
    instructions[3954] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 468 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 468, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3955] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 468 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 468, 'op': 'load'}
    instructions[3956] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 468 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 468, 'op': 'add'}
    instructions[3957] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 468 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 468, 'op': 'addl'}
    instructions[3958] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 468 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 468, 'op': 'load'}
    instructions[3959] = {5'd0, 4'd2, 4'd0, 16'd627};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 468 {'literal': 627, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 468, 'op': 'literal'}
    instructions[3960] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 468 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 468, 'op': 'store'}
    instructions[3961] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471, 'op': 'literal'}
    instructions[3962] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471, 'op': 'store'}
    instructions[3963] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471, 'op': 'addl'}
    instructions[3964] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471, 'op': 'addl'}
    instructions[3965] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471, 'op': 'addl'}
    instructions[3966] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471, 'op': 'load'}
    instructions[3967] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471, 'op': 'store'}
    instructions[3968] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471, 'op': 'addl'}
    instructions[3969] = {5'd0, 4'd8, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471 {'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471, 'op': 'literal'}
    instructions[3970] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471, 'op': 'store'}
    instructions[3971] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471, 'op': 'addl'}
    instructions[3972] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471, 'op': 'addl'}
    instructions[3973] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471, 'op': 'addl'}
    instructions[3974] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471, 'op': 'load'}
    instructions[3975] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3976] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471, 'op': 'load'}
    instructions[3977] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471, 'op': 'add'}
    instructions[3978] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3979] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471, 'op': 'load'}
    instructions[3980] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471, 'op': 'add'}
    instructions[3981] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471, 'op': 'addl'}
    instructions[3982] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471, 'op': 'load'}
    instructions[3983] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3984] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471, 'op': 'load'}
    instructions[3985] = {5'd22, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471, 'op': 'and'}
    instructions[3986] = {5'd0, 4'd2, 4'd0, 16'd586};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471 {'literal': 586, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471, 'op': 'literal'}
    instructions[3987] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 471, 'op': 'store'}
    instructions[3988] = {5'd0, 4'd8, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472 {'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472, 'op': 'literal'}
    instructions[3989] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472, 'op': 'store'}
    instructions[3990] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472, 'op': 'addl'}
    instructions[3991] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472, 'op': 'addl'}
    instructions[3992] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472, 'op': 'addl'}
    instructions[3993] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472, 'op': 'load'}
    instructions[3994] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472, 'op': 'store'}
    instructions[3995] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472, 'op': 'addl'}
    instructions[3996] = {5'd0, 4'd8, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472 {'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472, 'op': 'literal'}
    instructions[3997] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472, 'op': 'store'}
    instructions[3998] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472, 'op': 'addl'}
    instructions[3999] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472, 'op': 'addl'}
    instructions[4000] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472, 'op': 'addl'}
    instructions[4001] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472, 'op': 'load'}
    instructions[4002] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4003] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472, 'op': 'load'}
    instructions[4004] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472, 'op': 'add'}
    instructions[4005] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4006] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472, 'op': 'load'}
    instructions[4007] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472, 'op': 'add'}
    instructions[4008] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472, 'op': 'addl'}
    instructions[4009] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472, 'op': 'load'}
    instructions[4010] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4011] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472, 'op': 'load'}
    instructions[4012] = {5'd22, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472, 'op': 'and'}
    instructions[4013] = {5'd0, 4'd2, 4'd0, 16'd645};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472 {'literal': 645, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472, 'op': 'literal'}
    instructions[4014] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 472, 'op': 'store'}
    instructions[4015] = {5'd0, 4'd8, 4'd0, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473 {'literal': 4, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473, 'op': 'literal'}
    instructions[4016] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473, 'op': 'store'}
    instructions[4017] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473, 'op': 'addl'}
    instructions[4018] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473, 'op': 'addl'}
    instructions[4019] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473, 'op': 'addl'}
    instructions[4020] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473, 'op': 'load'}
    instructions[4021] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473, 'op': 'store'}
    instructions[4022] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473, 'op': 'addl'}
    instructions[4023] = {5'd0, 4'd8, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473 {'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473, 'op': 'literal'}
    instructions[4024] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473, 'op': 'store'}
    instructions[4025] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473, 'op': 'addl'}
    instructions[4026] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473, 'op': 'addl'}
    instructions[4027] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473, 'op': 'addl'}
    instructions[4028] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473, 'op': 'load'}
    instructions[4029] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4030] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473, 'op': 'load'}
    instructions[4031] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473, 'op': 'add'}
    instructions[4032] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4033] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473, 'op': 'load'}
    instructions[4034] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473, 'op': 'add'}
    instructions[4035] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473, 'op': 'addl'}
    instructions[4036] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473, 'op': 'load'}
    instructions[4037] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4038] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473, 'op': 'load'}
    instructions[4039] = {5'd22, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473, 'op': 'and'}
    instructions[4040] = {5'd0, 4'd2, 4'd0, 16'd587};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473 {'literal': 587, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473, 'op': 'literal'}
    instructions[4041] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 473, 'op': 'store'}
    instructions[4042] = {5'd0, 4'd8, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474 {'literal': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474, 'op': 'literal'}
    instructions[4043] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474, 'op': 'store'}
    instructions[4044] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474, 'op': 'addl'}
    instructions[4045] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474, 'op': 'addl'}
    instructions[4046] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474, 'op': 'addl'}
    instructions[4047] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474, 'op': 'load'}
    instructions[4048] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474, 'op': 'store'}
    instructions[4049] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474, 'op': 'addl'}
    instructions[4050] = {5'd0, 4'd8, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474 {'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474, 'op': 'literal'}
    instructions[4051] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474, 'op': 'store'}
    instructions[4052] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474, 'op': 'addl'}
    instructions[4053] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474, 'op': 'addl'}
    instructions[4054] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474, 'op': 'addl'}
    instructions[4055] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474, 'op': 'load'}
    instructions[4056] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4057] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474, 'op': 'load'}
    instructions[4058] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474, 'op': 'add'}
    instructions[4059] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4060] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474, 'op': 'load'}
    instructions[4061] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474, 'op': 'add'}
    instructions[4062] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474, 'op': 'addl'}
    instructions[4063] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474, 'op': 'load'}
    instructions[4064] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4065] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474, 'op': 'load'}
    instructions[4066] = {5'd22, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474, 'op': 'and'}
    instructions[4067] = {5'd0, 4'd2, 4'd0, 16'd25};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474 {'literal': 25, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474, 'op': 'literal'}
    instructions[4068] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 474, 'op': 'store'}
    instructions[4069] = {5'd0, 4'd8, 4'd0, 16'd16};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475 {'literal': 16, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475, 'op': 'literal'}
    instructions[4070] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475, 'op': 'store'}
    instructions[4071] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475, 'op': 'addl'}
    instructions[4072] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475, 'op': 'addl'}
    instructions[4073] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475, 'op': 'addl'}
    instructions[4074] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475, 'op': 'load'}
    instructions[4075] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475, 'op': 'store'}
    instructions[4076] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475, 'op': 'addl'}
    instructions[4077] = {5'd0, 4'd8, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475 {'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475, 'op': 'literal'}
    instructions[4078] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475, 'op': 'store'}
    instructions[4079] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475, 'op': 'addl'}
    instructions[4080] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475, 'op': 'addl'}
    instructions[4081] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475, 'op': 'addl'}
    instructions[4082] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475, 'op': 'load'}
    instructions[4083] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4084] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475, 'op': 'load'}
    instructions[4085] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475, 'op': 'add'}
    instructions[4086] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4087] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475, 'op': 'load'}
    instructions[4088] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475, 'op': 'add'}
    instructions[4089] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475, 'op': 'addl'}
    instructions[4090] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475, 'op': 'load'}
    instructions[4091] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4092] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475, 'op': 'load'}
    instructions[4093] = {5'd22, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475, 'op': 'and'}
    instructions[4094] = {5'd0, 4'd2, 4'd0, 16'd563};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475 {'literal': 563, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475, 'op': 'literal'}
    instructions[4095] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 475, 'op': 'store'}
    instructions[4096] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476, 'op': 'literal'}
    instructions[4097] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476, 'op': 'store'}
    instructions[4098] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476, 'op': 'addl'}
    instructions[4099] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476, 'op': 'addl'}
    instructions[4100] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476, 'op': 'addl'}
    instructions[4101] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476, 'op': 'load'}
    instructions[4102] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476, 'op': 'store'}
    instructions[4103] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476, 'op': 'addl'}
    instructions[4104] = {5'd0, 4'd8, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476 {'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476, 'op': 'literal'}
    instructions[4105] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476, 'op': 'store'}
    instructions[4106] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476, 'op': 'addl'}
    instructions[4107] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476, 'op': 'addl'}
    instructions[4108] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476, 'op': 'addl'}
    instructions[4109] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476, 'op': 'load'}
    instructions[4110] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4111] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476, 'op': 'load'}
    instructions[4112] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476, 'op': 'add'}
    instructions[4113] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4114] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476, 'op': 'load'}
    instructions[4115] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476, 'op': 'add'}
    instructions[4116] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476, 'op': 'addl'}
    instructions[4117] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476, 'op': 'load'}
    instructions[4118] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4119] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476, 'op': 'load'}
    instructions[4120] = {5'd22, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476, 'op': 'and'}
    instructions[4121] = {5'd0, 4'd2, 4'd0, 16'd542};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476 {'literal': 542, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476, 'op': 'literal'}
    instructions[4122] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 476, 'op': 'store'}
    instructions[4123] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 478 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 478, 'op': 'addl'}
    instructions[4124] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 478 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 478, 'op': 'addl'}
    instructions[4125] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 478 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 478, 'op': 'load'}
    instructions[4126] = {5'd0, 4'd2, 4'd0, 16'd646};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 478 {'literal': 646, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 478, 'op': 'literal'}
    instructions[4127] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 478 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 478, 'op': 'store'}
    instructions[4128] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 478 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 478, 'op': 'addl'}
    instructions[4129] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 478 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 478, 'op': 'addl'}
    instructions[4130] = {5'd16, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 478 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 478, 'op': 'return'}
    instructions[4131] = {5'd1, 4'd3, 4'd3, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 303 {'a': 3, 'literal': 10, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 303, 'op': 'addl'}
    instructions[4132] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 313 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 313, 'op': 'store'}
    instructions[4133] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 313 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 313, 'op': 'addl'}
    instructions[4134] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 313 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 313, 'op': 'store'}
    instructions[4135] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 313 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 313, 'op': 'addl'}
    instructions[4136] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 313 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 313, 'op': 'addl'}
    instructions[4137] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 313 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 313, 'op': 'addl'}
    instructions[4138] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 313 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 313, 'op': 'load'}
    instructions[4139] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 313 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 313, 'op': 'store'}
    instructions[4140] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 313 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 313, 'op': 'addl'}
    instructions[4141] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 313 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 313, 'op': 'addl'}
    instructions[4142] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 313 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 313, 'op': 'addl'}
    instructions[4143] = {5'd4, 4'd6, 4'd0, 16'd4654};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 313 {'z': 6, 'label': 4654, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 313, 'op': 'call'}
    instructions[4144] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 313 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 313, 'op': 'addl'}
    instructions[4145] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 313 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 313, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4146] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 313 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 313, 'op': 'load'}
    instructions[4147] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 313 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 313, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4148] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 313 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 313, 'op': 'load'}
    instructions[4149] = {5'd0, 4'd2, 4'd0, 16'd591};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 313 {'literal': 591, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 313, 'op': 'literal'}
    instructions[4150] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 313 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 313, 'op': 'load'}
    instructions[4151] = {5'd1, 4'd2, 4'd4, 16'd9};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 313 {'a': 4, 'literal': 9, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 313, 'op': 'addl'}
    instructions[4152] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 313 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 313, 'op': 'store'}
    instructions[4153] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 315 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 315, 'op': 'literal'}
    instructions[4154] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 315 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 315, 'op': 'store'}
    instructions[4155] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 315 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 315, 'op': 'addl'}
    instructions[4156] = {5'd1, 4'd8, 4'd4, 16'd9};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 315 {'a': 4, 'literal': 9, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 315, 'op': 'addl'}
    instructions[4157] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 315 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 315, 'op': 'addl'}
    instructions[4158] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 315 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 315, 'op': 'load'}
    instructions[4159] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 315 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 315, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4160] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 315 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 315, 'op': 'load'}
    instructions[4161] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 315 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 315, 'op': 'equal'}
    instructions[4162] = {5'd8, 4'd0, 4'd8, 16'd4170};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 315 {'a': 8, 'label': 4170, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 315, 'op': 'jmp_if_false'}
    instructions[4163] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 315 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 315, 'op': 'literal'}
    instructions[4164] = {5'd0, 4'd2, 4'd0, 16'd17};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 315 {'literal': 17, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 315, 'op': 'literal'}
    instructions[4165] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 315 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 315, 'op': 'store'}
    instructions[4166] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 315 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 315, 'op': 'addl'}
    instructions[4167] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 315 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 315, 'op': 'addl'}
    instructions[4168] = {5'd16, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 315 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 315, 'op': 'return'}
    instructions[4169] = {5'd10, 4'd0, 4'd0, 16'd4170};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 315 {'label': 4170, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 315, 'op': 'goto'}
    instructions[4170] = {5'd0, 4'd8, 4'd0, 16'd2048};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316 {'literal': 2048, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316, 'op': 'literal'}
    instructions[4171] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316, 'op': 'store'}
    instructions[4172] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316, 'op': 'addl'}
    instructions[4173] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316, 'op': 'addl'}
    instructions[4174] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316, 'op': 'addl'}
    instructions[4175] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316, 'op': 'load'}
    instructions[4176] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316, 'op': 'store'}
    instructions[4177] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316, 'op': 'addl'}
    instructions[4178] = {5'd0, 4'd8, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316 {'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316, 'op': 'literal'}
    instructions[4179] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4180] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316, 'op': 'load'}
    instructions[4181] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316, 'op': 'add'}
    instructions[4182] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316, 'op': 'addl'}
    instructions[4183] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316, 'op': 'load'}
    instructions[4184] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4185] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316, 'op': 'load'}
    instructions[4186] = {5'd13, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316, 'op': 'not_equal'}
    instructions[4187] = {5'd8, 4'd0, 4'd8, 16'd4195};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316 {'a': 8, 'label': 4195, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316, 'op': 'jmp_if_false'}
    instructions[4188] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316, 'op': 'literal'}
    instructions[4189] = {5'd0, 4'd2, 4'd0, 16'd17};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316 {'literal': 17, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316, 'op': 'literal'}
    instructions[4190] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316, 'op': 'store'}
    instructions[4191] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316, 'op': 'addl'}
    instructions[4192] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316, 'op': 'addl'}
    instructions[4193] = {5'd16, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316, 'op': 'return'}
    instructions[4194] = {5'd10, 4'd0, 4'd0, 16'd4195};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316 {'label': 4195, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 316, 'op': 'goto'}
    instructions[4195] = {5'd0, 4'd8, 4'd0, 16'd49320};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317 {'literal': 49320, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317, 'op': 'literal'}
    instructions[4196] = {5'd3, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317 {'a': 8, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317, 'op': 'literal_hi'}
    instructions[4197] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317, 'op': 'store'}
    instructions[4198] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317, 'op': 'addl'}
    instructions[4199] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317, 'op': 'addl'}
    instructions[4200] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317, 'op': 'addl'}
    instructions[4201] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317, 'op': 'load'}
    instructions[4202] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317, 'op': 'store'}
    instructions[4203] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317, 'op': 'addl'}
    instructions[4204] = {5'd0, 4'd8, 4'd0, 16'd15};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317 {'literal': 15, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317, 'op': 'literal'}
    instructions[4205] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4206] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317, 'op': 'load'}
    instructions[4207] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317, 'op': 'add'}
    instructions[4208] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317, 'op': 'addl'}
    instructions[4209] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317, 'op': 'load'}
    instructions[4210] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4211] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317, 'op': 'load'}
    instructions[4212] = {5'd13, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317, 'op': 'not_equal'}
    instructions[4213] = {5'd8, 4'd0, 4'd8, 16'd4221};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317 {'a': 8, 'label': 4221, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317, 'op': 'jmp_if_false'}
    instructions[4214] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317, 'op': 'literal'}
    instructions[4215] = {5'd0, 4'd2, 4'd0, 16'd17};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317 {'literal': 17, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317, 'op': 'literal'}
    instructions[4216] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317, 'op': 'store'}
    instructions[4217] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317, 'op': 'addl'}
    instructions[4218] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317, 'op': 'addl'}
    instructions[4219] = {5'd16, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317, 'op': 'return'}
    instructions[4220] = {5'd10, 4'd0, 4'd0, 16'd4221};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317 {'label': 4221, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 317, 'op': 'goto'}
    instructions[4221] = {5'd0, 4'd8, 4'd0, 16'd257};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318 {'literal': 257, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318, 'op': 'literal'}
    instructions[4222] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318, 'op': 'store'}
    instructions[4223] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318, 'op': 'addl'}
    instructions[4224] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318, 'op': 'addl'}
    instructions[4225] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318, 'op': 'addl'}
    instructions[4226] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318, 'op': 'load'}
    instructions[4227] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318, 'op': 'store'}
    instructions[4228] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318, 'op': 'addl'}
    instructions[4229] = {5'd0, 4'd8, 4'd0, 16'd16};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318 {'literal': 16, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318, 'op': 'literal'}
    instructions[4230] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4231] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318, 'op': 'load'}
    instructions[4232] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318, 'op': 'add'}
    instructions[4233] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318, 'op': 'addl'}
    instructions[4234] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318, 'op': 'load'}
    instructions[4235] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4236] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318, 'op': 'load'}
    instructions[4237] = {5'd13, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318, 'op': 'not_equal'}
    instructions[4238] = {5'd8, 4'd0, 4'd8, 16'd4246};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318 {'a': 8, 'label': 4246, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318, 'op': 'jmp_if_false'}
    instructions[4239] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318, 'op': 'literal'}
    instructions[4240] = {5'd0, 4'd2, 4'd0, 16'd17};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318 {'literal': 17, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318, 'op': 'literal'}
    instructions[4241] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318, 'op': 'store'}
    instructions[4242] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318, 'op': 'addl'}
    instructions[4243] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318, 'op': 'addl'}
    instructions[4244] = {5'd16, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318, 'op': 'return'}
    instructions[4245] = {5'd10, 4'd0, 4'd0, 16'd4246};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318 {'label': 4246, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 318, 'op': 'goto'}
    instructions[4246] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319, 'op': 'literal'}
    instructions[4247] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319, 'op': 'store'}
    instructions[4248] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319, 'op': 'addl'}
    instructions[4249] = {5'd0, 4'd8, 4'd0, 16'd255};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319 {'literal': 255, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319, 'op': 'literal'}
    instructions[4250] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319, 'op': 'store'}
    instructions[4251] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319, 'op': 'addl'}
    instructions[4252] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319, 'op': 'addl'}
    instructions[4253] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319, 'op': 'addl'}
    instructions[4254] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319, 'op': 'load'}
    instructions[4255] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319, 'op': 'store'}
    instructions[4256] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319, 'op': 'addl'}
    instructions[4257] = {5'd0, 4'd8, 4'd0, 16'd11};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319 {'literal': 11, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319, 'op': 'literal'}
    instructions[4258] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4259] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319, 'op': 'load'}
    instructions[4260] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319, 'op': 'add'}
    instructions[4261] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319, 'op': 'addl'}
    instructions[4262] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319, 'op': 'load'}
    instructions[4263] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4264] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319, 'op': 'load'}
    instructions[4265] = {5'd22, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319, 'op': 'and'}
    instructions[4266] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4267] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319, 'op': 'load'}
    instructions[4268] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319, 'op': 'equal'}
    instructions[4269] = {5'd8, 4'd0, 4'd8, 16'd4615};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319 {'a': 8, 'label': 4615, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319, 'op': 'jmp_if_false'}
    instructions[4270] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320, 'op': 'literal'}
    instructions[4271] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320, 'op': 'store'}
    instructions[4272] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320, 'op': 'addl'}
    instructions[4273] = {5'd0, 4'd8, 4'd0, 16'd15};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320 {'literal': 15, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320, 'op': 'literal'}
    instructions[4274] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320, 'op': 'store'}
    instructions[4275] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320, 'op': 'addl'}
    instructions[4276] = {5'd0, 4'd8, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320 {'literal': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320, 'op': 'literal'}
    instructions[4277] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320, 'op': 'store'}
    instructions[4278] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320, 'op': 'addl'}
    instructions[4279] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320, 'op': 'addl'}
    instructions[4280] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320, 'op': 'addl'}
    instructions[4281] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320, 'op': 'load'}
    instructions[4282] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320, 'op': 'store'}
    instructions[4283] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320, 'op': 'addl'}
    instructions[4284] = {5'd0, 4'd8, 4'd0, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320 {'literal': 7, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320, 'op': 'literal'}
    instructions[4285] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4286] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320, 'op': 'load'}
    instructions[4287] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320, 'op': 'add'}
    instructions[4288] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320, 'op': 'addl'}
    instructions[4289] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320, 'op': 'load'}
    instructions[4290] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4291] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320, 'op': 'load'}
    instructions[4292] = {5'd27, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320, 'op': 'shift_right'}
    instructions[4293] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4294] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320, 'op': 'load'}
    instructions[4295] = {5'd22, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320, 'op': 'and'}
    instructions[4296] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4297] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320, 'op': 'load'}
    instructions[4298] = {5'd28, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320, 'op': 'shift_left'}
    instructions[4299] = {5'd1, 4'd2, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320 {'a': 4, 'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320, 'op': 'addl'}
    instructions[4300] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 320, 'op': 'store'}
    instructions[4301] = {5'd0, 4'd8, 4'd0, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 321 {'literal': 7, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 321, 'op': 'literal'}
    instructions[4302] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 321 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 321, 'op': 'store'}
    instructions[4303] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 321 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 321, 'op': 'addl'}
    instructions[4304] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 321 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 321, 'op': 'addl'}
    instructions[4305] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 321 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 321, 'op': 'addl'}
    instructions[4306] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 321 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 321, 'op': 'load'}
    instructions[4307] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 321 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 321, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4308] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 321 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 321, 'op': 'load'}
    instructions[4309] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 321 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 321, 'op': 'add'}
    instructions[4310] = {5'd1, 4'd2, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 321 {'a': 4, 'literal': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 321, 'op': 'addl'}
    instructions[4311] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 321 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 321, 'op': 'store'}
    instructions[4312] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 322 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 322, 'op': 'addl'}
    instructions[4313] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 322 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 322, 'op': 'addl'}
    instructions[4314] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 322 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 322, 'op': 'load'}
    instructions[4315] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 322 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 322, 'op': 'store'}
    instructions[4316] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 322 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 322, 'op': 'addl'}
    instructions[4317] = {5'd0, 4'd8, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 322 {'literal': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 322, 'op': 'literal'}
    instructions[4318] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 322 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 322, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4319] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 322 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 322, 'op': 'load'}
    instructions[4320] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 322 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 322, 'op': 'add'}
    instructions[4321] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 322 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 322, 'op': 'addl'}
    instructions[4322] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 322 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 322, 'op': 'load'}
    instructions[4323] = {5'd1, 4'd2, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 322 {'a': 4, 'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 322, 'op': 'addl'}
    instructions[4324] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 322 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 322, 'op': 'store'}
    instructions[4325] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323, 'op': 'addl'}
    instructions[4326] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323, 'op': 'addl'}
    instructions[4327] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323, 'op': 'load'}
    instructions[4328] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323, 'op': 'store'}
    instructions[4329] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323, 'op': 'addl'}
    instructions[4330] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323, 'op': 'literal'}
    instructions[4331] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323, 'op': 'store'}
    instructions[4332] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323, 'op': 'addl'}
    instructions[4333] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323, 'op': 'literal'}
    instructions[4334] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323, 'op': 'store'}
    instructions[4335] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323, 'op': 'addl'}
    instructions[4336] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323, 'op': 'addl'}
    instructions[4337] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323, 'op': 'addl'}
    instructions[4338] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323, 'op': 'load'}
    instructions[4339] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4340] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323, 'op': 'load'}
    instructions[4341] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323, 'op': 'add'}
    instructions[4342] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4343] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323, 'op': 'load'}
    instructions[4344] = {5'd18, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323, 'op': 'unsigned_shift_right'}
    instructions[4345] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4346] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323, 'op': 'load'}
    instructions[4347] = {5'd9, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323, 'op': 'subtract'}
    instructions[4348] = {5'd1, 4'd2, 4'd4, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323 {'a': 4, 'literal': 4, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323, 'op': 'addl'}
    instructions[4349] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 323, 'op': 'store'}
    instructions[4350] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 324 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 324, 'op': 'literal'}
    instructions[4351] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 324 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 324, 'op': 'store'}
    instructions[4352] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 324 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 324, 'op': 'addl'}
    instructions[4353] = {5'd1, 4'd8, 4'd4, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 324 {'a': 4, 'literal': 4, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 324, 'op': 'addl'}
    instructions[4354] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 324 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 324, 'op': 'addl'}
    instructions[4355] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 324 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 324, 'op': 'load'}
    instructions[4356] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 324 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 324, 'op': 'store'}
    instructions[4357] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 324 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 324, 'op': 'addl'}
    instructions[4358] = {5'd1, 4'd8, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 324 {'a': 4, 'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 324, 'op': 'addl'}
    instructions[4359] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 324 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 324, 'op': 'addl'}
    instructions[4360] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 324 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 324, 'op': 'load'}
    instructions[4361] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 324 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 324, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4362] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 324 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 324, 'op': 'load'}
    instructions[4363] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 324 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 324, 'op': 'add'}
    instructions[4364] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 324 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 324, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4365] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 324 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 324, 'op': 'load'}
    instructions[4366] = {5'd9, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 324 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 324, 'op': 'subtract'}
    instructions[4367] = {5'd1, 4'd2, 4'd4, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 324 {'a': 4, 'literal': 8, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 324, 'op': 'addl'}
    instructions[4368] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 324 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 324, 'op': 'store'}
    instructions[4369] = {5'd0, 4'd8, 4'd0, 16'd2048};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 326 {'literal': 2048, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 326, 'op': 'literal'}
    instructions[4370] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 326 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 326, 'op': 'store'}
    instructions[4371] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 326 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 326, 'op': 'addl'}
    instructions[4372] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 326 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 326, 'op': 'addl'}
    instructions[4373] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 326 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 326, 'op': 'addl'}
    instructions[4374] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 326 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 326, 'op': 'load'}
    instructions[4375] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 326 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 326, 'op': 'store'}
    instructions[4376] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 326 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 326, 'op': 'addl'}
    instructions[4377] = {5'd1, 4'd8, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 326 {'a': 4, 'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 326, 'op': 'addl'}
    instructions[4378] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 326 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 326, 'op': 'addl'}
    instructions[4379] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 326 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 326, 'op': 'load'}
    instructions[4380] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 326 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 326, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4381] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 326 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 326, 'op': 'load'}
    instructions[4382] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 326 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 326, 'op': 'add'}
    instructions[4383] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 326 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 326, 'op': 'addl'}
    instructions[4384] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 326 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 326, 'op': 'load'}
    instructions[4385] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 326 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 326, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4386] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 326 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 326, 'op': 'load'}
    instructions[4387] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 326 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 326, 'op': 'equal'}
    instructions[4388] = {5'd8, 4'd0, 4'd8, 16'd4608};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 326 {'a': 8, 'label': 4608, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 326, 'op': 'jmp_if_false'}
    instructions[4389] = {5'd0, 4'd8, 4'd0, 16'd19};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 329 {'literal': 19, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 329, 'op': 'literal'}
    instructions[4390] = {5'd1, 4'd2, 4'd4, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 329 {'a': 4, 'literal': 7, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 329, 'op': 'addl'}
    instructions[4391] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 329 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 329, 'op': 'store'}
    instructions[4392] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 330 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 330, 'op': 'store'}
    instructions[4393] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 330 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 330, 'op': 'addl'}
    instructions[4394] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 330 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 330, 'op': 'store'}
    instructions[4395] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 330 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 330, 'op': 'addl'}
    instructions[4396] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 330 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 330, 'op': 'addl'}
    instructions[4397] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 330 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 330, 'op': 'addl'}
    instructions[4398] = {5'd4, 4'd6, 4'd0, 16'd1952};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 330 {'z': 6, 'label': 1952, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 330, 'op': 'call'}
    instructions[4399] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 330 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 330, 'op': 'addl'}
    instructions[4400] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 330 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 330, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4401] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 330 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 330, 'op': 'load'}
    instructions[4402] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 330 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 330, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4403] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 330 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 330, 'op': 'load'}
    instructions[4404] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 330 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 330, 'op': 'addl'}
    instructions[4405] = {5'd0, 4'd8, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331 {'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331, 'op': 'literal'}
    instructions[4406] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331, 'op': 'store'}
    instructions[4407] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331, 'op': 'addl'}
    instructions[4408] = {5'd1, 4'd8, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331 {'a': 4, 'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331, 'op': 'addl'}
    instructions[4409] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331, 'op': 'addl'}
    instructions[4410] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331, 'op': 'load'}
    instructions[4411] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4412] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331, 'op': 'load'}
    instructions[4413] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331, 'op': 'add'}
    instructions[4414] = {5'd1, 4'd2, 4'd4, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331 {'a': 4, 'literal': 6, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331, 'op': 'addl'}
    instructions[4415] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331, 'op': 'store'}
    instructions[4416] = {5'd1, 4'd8, 4'd4, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331 {'a': 4, 'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331, 'op': 'addl'}
    instructions[4417] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331, 'op': 'addl'}
    instructions[4418] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331, 'op': 'load'}
    instructions[4419] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331, 'op': 'store'}
    instructions[4420] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331, 'op': 'addl'}
    instructions[4421] = {5'd1, 4'd8, 4'd4, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331 {'a': 4, 'literal': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331, 'op': 'addl'}
    instructions[4422] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331, 'op': 'addl'}
    instructions[4423] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331, 'op': 'load'}
    instructions[4424] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4425] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331, 'op': 'load'}
    instructions[4426] = {5'd24, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331, 'op': 'unsigned_greater_equal'}
    instructions[4427] = {5'd8, 4'd0, 4'd8, 16'd4516};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331 {'a': 8, 'label': 4516, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331, 'op': 'jmp_if_false'}
    instructions[4428] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 332 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 332, 'op': 'addl'}
    instructions[4429] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 332 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 332, 'op': 'addl'}
    instructions[4430] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 332 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 332, 'op': 'load'}
    instructions[4431] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 332 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 332, 'op': 'store'}
    instructions[4432] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 332 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 332, 'op': 'addl'}
    instructions[4433] = {5'd1, 4'd8, 4'd4, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 332 {'a': 4, 'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 332, 'op': 'addl'}
    instructions[4434] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 332 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 332, 'op': 'addl'}
    instructions[4435] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 332 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 332, 'op': 'load'}
    instructions[4436] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 332 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 332, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4437] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 332 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 332, 'op': 'load'}
    instructions[4438] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 332 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 332, 'op': 'add'}
    instructions[4439] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 332 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 332, 'op': 'addl'}
    instructions[4440] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 332 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 332, 'op': 'load'}
    instructions[4441] = {5'd1, 4'd2, 4'd4, 16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 332 {'a': 4, 'literal': 5, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 332, 'op': 'addl'}
    instructions[4442] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 332 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 332, 'op': 'store'}
    instructions[4443] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 333 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 333, 'op': 'store'}
    instructions[4444] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 333 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 333, 'op': 'addl'}
    instructions[4445] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 333 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 333, 'op': 'store'}
    instructions[4446] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 333 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 333, 'op': 'addl'}
    instructions[4447] = {5'd1, 4'd8, 4'd4, 16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 333 {'a': 4, 'literal': 5, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 333, 'op': 'addl'}
    instructions[4448] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 333 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 333, 'op': 'addl'}
    instructions[4449] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 333 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 333, 'op': 'load'}
    instructions[4450] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 333 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 333, 'op': 'store'}
    instructions[4451] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 333 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 333, 'op': 'addl'}
    instructions[4452] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 333 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 333, 'op': 'addl'}
    instructions[4453] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 333 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 333, 'op': 'addl'}
    instructions[4454] = {5'd4, 4'd6, 4'd0, 16'd1962};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 333 {'z': 6, 'label': 1962, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 333, 'op': 'call'}
    instructions[4455] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 333 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 333, 'op': 'addl'}
    instructions[4456] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 333 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 333, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4457] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 333 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 333, 'op': 'load'}
    instructions[4458] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 333 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 333, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4459] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 333 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 333, 'op': 'load'}
    instructions[4460] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 333 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 333, 'op': 'addl'}
    instructions[4461] = {5'd1, 4'd8, 4'd4, 16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 334 {'a': 4, 'literal': 5, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 334, 'op': 'addl'}
    instructions[4462] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 334 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 334, 'op': 'addl'}
    instructions[4463] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 334 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 334, 'op': 'load'}
    instructions[4464] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 334 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 334, 'op': 'store'}
    instructions[4465] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 334 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 334, 'op': 'addl'}
    instructions[4466] = {5'd0, 4'd8, 4'd0, 16'd27};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 334 {'literal': 27, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 334, 'op': 'literal'}
    instructions[4467] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 334 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 334, 'op': 'store'}
    instructions[4468] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 334 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 334, 'op': 'addl'}
    instructions[4469] = {5'd1, 4'd8, 4'd4, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 334 {'a': 4, 'literal': 7, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 334, 'op': 'addl'}
    instructions[4470] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 334 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 334, 'op': 'addl'}
    instructions[4471] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 334 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 334, 'op': 'load'}
    instructions[4472] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 334 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 334, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4473] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 334 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 334, 'op': 'load'}
    instructions[4474] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 334 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 334, 'op': 'add'}
    instructions[4475] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 334 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 334, 'op': 'addl'}
    instructions[4476] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 334 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 334, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4477] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 334 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 334, 'op': 'load'}
    instructions[4478] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 334 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 334, 'op': 'store'}
    instructions[4479] = {5'd1, 4'd8, 4'd4, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 335 {'a': 4, 'literal': 7, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 335, 'op': 'addl'}
    instructions[4480] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 335 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 335, 'op': 'addl'}
    instructions[4481] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 335 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 335, 'op': 'load'}
    instructions[4482] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 335 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 335, 'op': 'store'}
    instructions[4483] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 335 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 335, 'op': 'addl'}
    instructions[4484] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 335 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 335, 'op': 'literal'}
    instructions[4485] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 335 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 335, 'op': 'store'}
    instructions[4486] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 335 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 335, 'op': 'addl'}
    instructions[4487] = {5'd1, 4'd8, 4'd4, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 335 {'a': 4, 'literal': 7, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 335, 'op': 'addl'}
    instructions[4488] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 335 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 335, 'op': 'addl'}
    instructions[4489] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 335 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 335, 'op': 'load'}
    instructions[4490] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 335 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 335, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4491] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 335 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 335, 'op': 'load'}
    instructions[4492] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 335 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 335, 'op': 'add'}
    instructions[4493] = {5'd1, 4'd2, 4'd4, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 335 {'a': 4, 'literal': 7, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 335, 'op': 'addl'}
    instructions[4494] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 335 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 335, 'op': 'store'}
    instructions[4495] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 335 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 335, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4496] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 335 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 335, 'op': 'load'}
    instructions[4497] = {5'd1, 4'd8, 4'd4, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331 {'a': 4, 'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331, 'op': 'addl'}
    instructions[4498] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331, 'op': 'addl'}
    instructions[4499] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331, 'op': 'load'}
    instructions[4500] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331, 'op': 'store'}
    instructions[4501] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331, 'op': 'addl'}
    instructions[4502] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331, 'op': 'literal'}
    instructions[4503] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331, 'op': 'store'}
    instructions[4504] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331, 'op': 'addl'}
    instructions[4505] = {5'd1, 4'd8, 4'd4, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331 {'a': 4, 'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331, 'op': 'addl'}
    instructions[4506] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331, 'op': 'addl'}
    instructions[4507] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331, 'op': 'load'}
    instructions[4508] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4509] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331, 'op': 'load'}
    instructions[4510] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331, 'op': 'add'}
    instructions[4511] = {5'd1, 4'd2, 4'd4, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331 {'a': 4, 'literal': 6, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331, 'op': 'addl'}
    instructions[4512] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331, 'op': 'store'}
    instructions[4513] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4514] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331, 'op': 'load'}
    instructions[4515] = {5'd10, 4'd0, 4'd0, 16'd4416};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331 {'label': 4416, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 331, 'op': 'goto'}
    instructions[4516] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 337 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 337, 'op': 'literal'}
    instructions[4517] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 337 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 337, 'op': 'store'}
    instructions[4518] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 337 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 337, 'op': 'addl'}
    instructions[4519] = {5'd0, 4'd8, 4'd0, 16'd27};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 337 {'literal': 27, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 337, 'op': 'literal'}
    instructions[4520] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 337 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 337, 'op': 'store'}
    instructions[4521] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 337 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 337, 'op': 'addl'}
    instructions[4522] = {5'd0, 4'd8, 4'd0, 16'd17};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 337 {'literal': 17, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 337, 'op': 'literal'}
    instructions[4523] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 337 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 337, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4524] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 337 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 337, 'op': 'load'}
    instructions[4525] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 337 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 337, 'op': 'add'}
    instructions[4526] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 337 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 337, 'op': 'addl'}
    instructions[4527] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 337 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 337, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4528] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 337 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 337, 'op': 'load'}
    instructions[4529] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 337 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 337, 'op': 'store'}
    instructions[4530] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338, 'op': 'store'}
    instructions[4531] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338, 'op': 'addl'}
    instructions[4532] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338, 'op': 'store'}
    instructions[4533] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338, 'op': 'addl'}
    instructions[4534] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338, 'op': 'addl'}
    instructions[4535] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338, 'op': 'addl'}
    instructions[4536] = {5'd4, 4'd6, 4'd0, 16'd2053};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338 {'z': 6, 'label': 2053, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338, 'op': 'call'}
    instructions[4537] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338, 'op': 'addl'}
    instructions[4538] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4539] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338, 'op': 'load'}
    instructions[4540] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4541] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338, 'op': 'load'}
    instructions[4542] = {5'd0, 4'd2, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338 {'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338, 'op': 'literal'}
    instructions[4543] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338, 'op': 'load'}
    instructions[4544] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338, 'op': 'store'}
    instructions[4545] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338, 'op': 'addl'}
    instructions[4546] = {5'd0, 4'd8, 4'd0, 16'd27};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338 {'literal': 27, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338, 'op': 'literal'}
    instructions[4547] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338, 'op': 'store'}
    instructions[4548] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338, 'op': 'addl'}
    instructions[4549] = {5'd0, 4'd8, 4'd0, 16'd18};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338 {'literal': 18, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338, 'op': 'literal'}
    instructions[4550] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4551] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338, 'op': 'load'}
    instructions[4552] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338, 'op': 'add'}
    instructions[4553] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338, 'op': 'addl'}
    instructions[4554] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4555] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338, 'op': 'load'}
    instructions[4556] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 338, 'op': 'store'}
    instructions[4557] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 341 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 341, 'op': 'store'}
    instructions[4558] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 341 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 341, 'op': 'addl'}
    instructions[4559] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 341 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 341, 'op': 'store'}
    instructions[4560] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 341 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 341, 'op': 'addl'}
    instructions[4561] = {5'd0, 4'd8, 4'd0, 16'd27};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 342 {'literal': 27, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 342, 'op': 'literal'}
    instructions[4562] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 341 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 341, 'op': 'store'}
    instructions[4563] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 341 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 341, 'op': 'addl'}
    instructions[4564] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 343 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 343, 'op': 'addl'}
    instructions[4565] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 343 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 343, 'op': 'addl'}
    instructions[4566] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 343 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 343, 'op': 'load'}
    instructions[4567] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 341 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 341, 'op': 'store'}
    instructions[4568] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 341 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 341, 'op': 'addl'}
    instructions[4569] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 344 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 344, 'op': 'literal'}
    instructions[4570] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 341 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 341, 'op': 'store'}
    instructions[4571] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 341 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 341, 'op': 'addl'}
    instructions[4572] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 345 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 345, 'op': 'addl'}
    instructions[4573] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 345 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 345, 'op': 'addl'}
    instructions[4574] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 345 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 345, 'op': 'load'}
    instructions[4575] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 345 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 345, 'op': 'store'}
    instructions[4576] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 345 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 345, 'op': 'addl'}
    instructions[4577] = {5'd0, 4'd8, 4'd0, 16'd13};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 345 {'literal': 13, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 345, 'op': 'literal'}
    instructions[4578] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 345 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 345, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4579] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 345 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 345, 'op': 'load'}
    instructions[4580] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 345 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 345, 'op': 'add'}
    instructions[4581] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 345 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 345, 'op': 'addl'}
    instructions[4582] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 345 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 345, 'op': 'load'}
    instructions[4583] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 341 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 341, 'op': 'store'}
    instructions[4584] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 341 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 341, 'op': 'addl'}
    instructions[4585] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 346 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 346, 'op': 'addl'}
    instructions[4586] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 346 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 346, 'op': 'addl'}
    instructions[4587] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 346 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 346, 'op': 'load'}
    instructions[4588] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 347 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 347, 'op': 'store'}
    instructions[4589] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 347 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 347, 'op': 'addl'}
    instructions[4590] = {5'd0, 4'd8, 4'd0, 16'd14};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 346 {'literal': 14, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 346, 'op': 'literal'}
    instructions[4591] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 347 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 347, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4592] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 347 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 347, 'op': 'load'}
    instructions[4593] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 347 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 347, 'op': 'add'}
    instructions[4594] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 347 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 347, 'op': 'addl'}
    instructions[4595] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 347 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 347, 'op': 'load'}
    instructions[4596] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 341 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 341, 'op': 'store'}
    instructions[4597] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 341 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 341, 'op': 'addl'}
    instructions[4598] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 341 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 341, 'op': 'addl'}
    instructions[4599] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 341 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 341, 'op': 'addl'}
    instructions[4600] = {5'd4, 4'd6, 4'd0, 16'd2066};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 341 {'z': 6, 'label': 2066, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 341, 'op': 'call'}
    instructions[4601] = {5'd1, 4'd3, 4'd3, -16'd5};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 341 {'a': 3, 'literal': -5, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 341, 'op': 'addl'}
    instructions[4602] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 341 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 341, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4603] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 341 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 341, 'op': 'load'}
    instructions[4604] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 341 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 341, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4605] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 341 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 341, 'op': 'load'}
    instructions[4606] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 341 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 341, 'op': 'addl'}
    instructions[4607] = {5'd10, 4'd0, 4'd0, 16'd4608};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 326 {'label': 4608, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 326, 'op': 'goto'}
    instructions[4608] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 349 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 349, 'op': 'literal'}
    instructions[4609] = {5'd0, 4'd2, 4'd0, 16'd17};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 349 {'literal': 17, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 349, 'op': 'literal'}
    instructions[4610] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 349 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 349, 'op': 'store'}
    instructions[4611] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 349 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 349, 'op': 'addl'}
    instructions[4612] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 349 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 349, 'op': 'addl'}
    instructions[4613] = {5'd16, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 349 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 349, 'op': 'return'}
    instructions[4614] = {5'd10, 4'd0, 4'd0, 16'd4615};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319 {'label': 4615, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 319, 'op': 'goto'}
    instructions[4615] = {5'd0, 4'd8, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352 {'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352, 'op': 'literal'}
    instructions[4616] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352, 'op': 'store'}
    instructions[4617] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352, 'op': 'addl'}
    instructions[4618] = {5'd0, 4'd8, 4'd0, 16'd255};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352 {'literal': 255, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352, 'op': 'literal'}
    instructions[4619] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352, 'op': 'store'}
    instructions[4620] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352, 'op': 'addl'}
    instructions[4621] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352, 'op': 'addl'}
    instructions[4622] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352, 'op': 'addl'}
    instructions[4623] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352, 'op': 'load'}
    instructions[4624] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352, 'op': 'store'}
    instructions[4625] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352, 'op': 'addl'}
    instructions[4626] = {5'd0, 4'd8, 4'd0, 16'd11};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352 {'literal': 11, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352, 'op': 'literal'}
    instructions[4627] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4628] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352, 'op': 'load'}
    instructions[4629] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352, 'op': 'add'}
    instructions[4630] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352, 'op': 'addl'}
    instructions[4631] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352, 'op': 'load'}
    instructions[4632] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4633] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352, 'op': 'load'}
    instructions[4634] = {5'd22, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352, 'op': 'and'}
    instructions[4635] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4636] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352, 'op': 'load'}
    instructions[4637] = {5'd13, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352, 'op': 'not_equal'}
    instructions[4638] = {5'd8, 4'd0, 4'd8, 16'd4646};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352 {'a': 8, 'label': 4646, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352, 'op': 'jmp_if_false'}
    instructions[4639] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352, 'op': 'literal'}
    instructions[4640] = {5'd0, 4'd2, 4'd0, 16'd17};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352 {'literal': 17, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352, 'op': 'literal'}
    instructions[4641] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352, 'op': 'store'}
    instructions[4642] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352, 'op': 'addl'}
    instructions[4643] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352, 'op': 'addl'}
    instructions[4644] = {5'd16, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352, 'op': 'return'}
    instructions[4645] = {5'd10, 4'd0, 4'd0, 16'd4646};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352 {'label': 4646, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 352, 'op': 'goto'}
    instructions[4646] = {5'd1, 4'd8, 4'd4, 16'd9};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 353 {'a': 4, 'literal': 9, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 353, 'op': 'addl'}
    instructions[4647] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 353 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 353, 'op': 'addl'}
    instructions[4648] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 353 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 353, 'op': 'load'}
    instructions[4649] = {5'd0, 4'd2, 4'd0, 16'd17};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 353 {'literal': 17, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 353, 'op': 'literal'}
    instructions[4650] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 353 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 353, 'op': 'store'}
    instructions[4651] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 353 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 353, 'op': 'addl'}
    instructions[4652] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 353 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 353, 'op': 'addl'}
    instructions[4653] = {5'd16, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 353 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 353, 'op': 'return'}
    instructions[4654] = {5'd1, 4'd3, 4'd3, 16'd9};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 132 {'a': 3, 'literal': 9, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 132, 'op': 'addl'}
    instructions[4655] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137, 'op': 'literal'}
    instructions[4656] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137, 'op': 'store'}
    instructions[4657] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137, 'op': 'addl'}
    instructions[4658] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137, 'op': 'store'}
    instructions[4659] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137, 'op': 'addl'}
    instructions[4660] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137, 'op': 'store'}
    instructions[4661] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137, 'op': 'addl'}
    instructions[4662] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137, 'op': 'addl'}
    instructions[4663] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137, 'op': 'addl'}
    instructions[4664] = {5'd4, 4'd6, 4'd0, 16'd5286};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137 {'z': 6, 'label': 5286, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137, 'op': 'call'}
    instructions[4665] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137, 'op': 'addl'}
    instructions[4666] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4667] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137, 'op': 'load'}
    instructions[4668] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4669] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137, 'op': 'load'}
    instructions[4670] = {5'd0, 4'd2, 4'd0, 16'd26};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137 {'literal': 26, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137, 'op': 'literal'}
    instructions[4671] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137, 'op': 'load'}
    instructions[4672] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4673] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137, 'op': 'load'}
    instructions[4674] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137, 'op': 'equal'}
    instructions[4675] = {5'd8, 4'd0, 4'd8, 16'd4683};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137 {'a': 8, 'label': 4683, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137, 'op': 'jmp_if_false'}
    instructions[4676] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137, 'op': 'literal'}
    instructions[4677] = {5'd0, 4'd2, 4'd0, 16'd591};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137 {'literal': 591, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137, 'op': 'literal'}
    instructions[4678] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137, 'op': 'store'}
    instructions[4679] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137, 'op': 'addl'}
    instructions[4680] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137, 'op': 'addl'}
    instructions[4681] = {5'd16, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137, 'op': 'return'}
    instructions[4682] = {5'd10, 4'd0, 4'd0, 16'd4683};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137 {'label': 4683, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 137, 'op': 'goto'}
    instructions[4683] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 139 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 139, 'op': 'store'}
    instructions[4684] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 139 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 139, 'op': 'addl'}
    instructions[4685] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 139 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 139, 'op': 'store'}
    instructions[4686] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 139 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 139, 'op': 'addl'}
    instructions[4687] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 139 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 139, 'op': 'addl'}
    instructions[4688] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 139 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 139, 'op': 'addl'}
    instructions[4689] = {5'd4, 4'd6, 4'd0, 16'd3315};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 139 {'z': 6, 'label': 3315, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 139, 'op': 'call'}
    instructions[4690] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 139 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 139, 'op': 'addl'}
    instructions[4691] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 139 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 139, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4692] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 139 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 139, 'op': 'load'}
    instructions[4693] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 139 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 139, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4694] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 139 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 139, 'op': 'load'}
    instructions[4695] = {5'd0, 4'd2, 4'd0, 16'd540};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 139 {'literal': 540, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 139, 'op': 'literal'}
    instructions[4696] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 139 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 139, 'op': 'load'}
    instructions[4697] = {5'd1, 4'd2, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 139 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 139, 'op': 'addl'}
    instructions[4698] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 139 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 139, 'op': 'store'}
    instructions[4699] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 140 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 140, 'op': 'literal'}
    instructions[4700] = {5'd1, 4'd2, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 140 {'a': 4, 'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 140, 'op': 'addl'}
    instructions[4701] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 140 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 140, 'op': 'store'}
    instructions[4702] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141, 'op': 'literal'}
    instructions[4703] = {5'd1, 4'd2, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141 {'a': 4, 'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141, 'op': 'addl'}
    instructions[4704] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141, 'op': 'store'}
    instructions[4705] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141, 'op': 'addl'}
    instructions[4706] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141, 'op': 'addl'}
    instructions[4707] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141, 'op': 'load'}
    instructions[4708] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141, 'op': 'store'}
    instructions[4709] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141, 'op': 'addl'}
    instructions[4710] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141, 'op': 'addl'}
    instructions[4711] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141, 'op': 'addl'}
    instructions[4712] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141, 'op': 'load'}
    instructions[4713] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4714] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141, 'op': 'load'}
    instructions[4715] = {5'd19, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141, 'op': 'unsigned_greater'}
    instructions[4716] = {5'd8, 4'd0, 4'd8, 16'd4778};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141 {'a': 8, 'label': 4778, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141, 'op': 'jmp_if_false'}
    instructions[4717] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142, 'op': 'store'}
    instructions[4718] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142, 'op': 'addl'}
    instructions[4719] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142, 'op': 'store'}
    instructions[4720] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142, 'op': 'addl'}
    instructions[4721] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142, 'op': 'addl'}
    instructions[4722] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142, 'op': 'addl'}
    instructions[4723] = {5'd4, 4'd6, 4'd0, 16'd3315};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142 {'z': 6, 'label': 3315, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142, 'op': 'call'}
    instructions[4724] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142, 'op': 'addl'}
    instructions[4725] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4726] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142, 'op': 'load'}
    instructions[4727] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4728] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142, 'op': 'load'}
    instructions[4729] = {5'd0, 4'd2, 4'd0, 16'd540};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142 {'literal': 540, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142, 'op': 'literal'}
    instructions[4730] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142, 'op': 'load'}
    instructions[4731] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142, 'op': 'store'}
    instructions[4732] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142, 'op': 'addl'}
    instructions[4733] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142, 'op': 'addl'}
    instructions[4734] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142, 'op': 'addl'}
    instructions[4735] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142, 'op': 'load'}
    instructions[4736] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142, 'op': 'store'}
    instructions[4737] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142, 'op': 'addl'}
    instructions[4738] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142, 'op': 'addl'}
    instructions[4739] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142, 'op': 'addl'}
    instructions[4740] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142, 'op': 'load'}
    instructions[4741] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4742] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142, 'op': 'load'}
    instructions[4743] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142, 'op': 'add'}
    instructions[4744] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142, 'op': 'addl'}
    instructions[4745] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4746] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142, 'op': 'load'}
    instructions[4747] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 142, 'op': 'store'}
    instructions[4748] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 143 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 143, 'op': 'addl'}
    instructions[4749] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 143 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 143, 'op': 'addl'}
    instructions[4750] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 143 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 143, 'op': 'load'}
    instructions[4751] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 143 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 143, 'op': 'store'}
    instructions[4752] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 143 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 143, 'op': 'addl'}
    instructions[4753] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 143 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 143, 'op': 'literal'}
    instructions[4754] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 143 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 143, 'op': 'store'}
    instructions[4755] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 143 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 143, 'op': 'addl'}
    instructions[4756] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 143 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 143, 'op': 'addl'}
    instructions[4757] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 143 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 143, 'op': 'addl'}
    instructions[4758] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 143 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 143, 'op': 'load'}
    instructions[4759] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 143 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 143, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4760] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 143 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 143, 'op': 'load'}
    instructions[4761] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 143 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 143, 'op': 'add'}
    instructions[4762] = {5'd1, 4'd2, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 143 {'a': 4, 'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 143, 'op': 'addl'}
    instructions[4763] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 143 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 143, 'op': 'store'}
    instructions[4764] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 143 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 143, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4765] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 143 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 143, 'op': 'load'}
    instructions[4766] = {5'd0, 4'd8, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141 {'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141, 'op': 'literal'}
    instructions[4767] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141, 'op': 'store'}
    instructions[4768] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141, 'op': 'addl'}
    instructions[4769] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141, 'op': 'addl'}
    instructions[4770] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141, 'op': 'addl'}
    instructions[4771] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141, 'op': 'load'}
    instructions[4772] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4773] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141, 'op': 'load'}
    instructions[4774] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141, 'op': 'add'}
    instructions[4775] = {5'd1, 4'd2, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141 {'a': 4, 'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141, 'op': 'addl'}
    instructions[4776] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141, 'op': 'store'}
    instructions[4777] = {5'd10, 4'd0, 4'd0, 16'd4705};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141 {'label': 4705, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 141, 'op': 'goto'}
    instructions[4778] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147, 'op': 'literal'}
    instructions[4779] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147, 'op': 'store'}
    instructions[4780] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147, 'op': 'addl'}
    instructions[4781] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147, 'op': 'addl'}
    instructions[4782] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147, 'op': 'addl'}
    instructions[4783] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147, 'op': 'load'}
    instructions[4784] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147, 'op': 'store'}
    instructions[4785] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147, 'op': 'addl'}
    instructions[4786] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147, 'op': 'literal'}
    instructions[4787] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4788] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147, 'op': 'load'}
    instructions[4789] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147, 'op': 'add'}
    instructions[4790] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147, 'op': 'addl'}
    instructions[4791] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147, 'op': 'load'}
    instructions[4792] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4793] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147, 'op': 'load'}
    instructions[4794] = {5'd13, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147, 'op': 'not_equal'}
    instructions[4795] = {5'd8, 4'd0, 4'd8, 16'd4814};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147 {'a': 8, 'label': 4814, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147, 'op': 'jmp_if_false'}
    instructions[4796] = {5'd0, 4'd8, 4'd0, 16'd65535};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147 {'literal': 65535, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147, 'op': 'literal'}
    instructions[4797] = {5'd3, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147 {'a': 8, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147, 'op': 'literal_hi'}
    instructions[4798] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147, 'op': 'store'}
    instructions[4799] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147, 'op': 'addl'}
    instructions[4800] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147, 'op': 'addl'}
    instructions[4801] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147, 'op': 'addl'}
    instructions[4802] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147, 'op': 'load'}
    instructions[4803] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147, 'op': 'store'}
    instructions[4804] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147, 'op': 'addl'}
    instructions[4805] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147, 'op': 'literal'}
    instructions[4806] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4807] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147, 'op': 'load'}
    instructions[4808] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147, 'op': 'add'}
    instructions[4809] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147, 'op': 'addl'}
    instructions[4810] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147, 'op': 'load'}
    instructions[4811] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4812] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147, 'op': 'load'}
    instructions[4813] = {5'd13, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147, 'op': 'not_equal'}
    instructions[4814] = {5'd8, 4'd0, 4'd8, 16'd4822};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147 {'a': 8, 'label': 4822, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147, 'op': 'jmp_if_false'}
    instructions[4815] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147, 'op': 'literal'}
    instructions[4816] = {5'd0, 4'd2, 4'd0, 16'd591};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147 {'literal': 591, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147, 'op': 'literal'}
    instructions[4817] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147, 'op': 'store'}
    instructions[4818] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147, 'op': 'addl'}
    instructions[4819] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147, 'op': 'addl'}
    instructions[4820] = {5'd16, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147, 'op': 'return'}
    instructions[4821] = {5'd10, 4'd0, 4'd0, 16'd4822};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147 {'label': 4822, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 147, 'op': 'goto'}
    instructions[4822] = {5'd0, 4'd8, 4'd0, 16'd515};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148 {'literal': 515, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148, 'op': 'literal'}
    instructions[4823] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148, 'op': 'store'}
    instructions[4824] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148, 'op': 'addl'}
    instructions[4825] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148, 'op': 'addl'}
    instructions[4826] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148, 'op': 'addl'}
    instructions[4827] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148, 'op': 'load'}
    instructions[4828] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148, 'op': 'store'}
    instructions[4829] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148, 'op': 'addl'}
    instructions[4830] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148, 'op': 'literal'}
    instructions[4831] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4832] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148, 'op': 'load'}
    instructions[4833] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148, 'op': 'add'}
    instructions[4834] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148, 'op': 'addl'}
    instructions[4835] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148, 'op': 'load'}
    instructions[4836] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4837] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148, 'op': 'load'}
    instructions[4838] = {5'd13, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148, 'op': 'not_equal'}
    instructions[4839] = {5'd8, 4'd0, 4'd8, 16'd4858};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148 {'a': 8, 'label': 4858, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148, 'op': 'jmp_if_false'}
    instructions[4840] = {5'd0, 4'd8, 4'd0, 16'd65535};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148 {'literal': 65535, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148, 'op': 'literal'}
    instructions[4841] = {5'd3, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148 {'a': 8, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148, 'op': 'literal_hi'}
    instructions[4842] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148, 'op': 'store'}
    instructions[4843] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148, 'op': 'addl'}
    instructions[4844] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148, 'op': 'addl'}
    instructions[4845] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148, 'op': 'addl'}
    instructions[4846] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148, 'op': 'load'}
    instructions[4847] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148, 'op': 'store'}
    instructions[4848] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148, 'op': 'addl'}
    instructions[4849] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148, 'op': 'literal'}
    instructions[4850] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4851] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148, 'op': 'load'}
    instructions[4852] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148, 'op': 'add'}
    instructions[4853] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148, 'op': 'addl'}
    instructions[4854] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148, 'op': 'load'}
    instructions[4855] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4856] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148, 'op': 'load'}
    instructions[4857] = {5'd13, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148, 'op': 'not_equal'}
    instructions[4858] = {5'd8, 4'd0, 4'd8, 16'd4866};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148 {'a': 8, 'label': 4866, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148, 'op': 'jmp_if_false'}
    instructions[4859] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148, 'op': 'literal'}
    instructions[4860] = {5'd0, 4'd2, 4'd0, 16'd591};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148 {'literal': 591, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148, 'op': 'literal'}
    instructions[4861] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148, 'op': 'store'}
    instructions[4862] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148, 'op': 'addl'}
    instructions[4863] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148, 'op': 'addl'}
    instructions[4864] = {5'd16, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148, 'op': 'return'}
    instructions[4865] = {5'd10, 4'd0, 4'd0, 16'd4866};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148 {'label': 4866, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 148, 'op': 'goto'}
    instructions[4866] = {5'd0, 4'd8, 4'd0, 16'd1029};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149 {'literal': 1029, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149, 'op': 'literal'}
    instructions[4867] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149, 'op': 'store'}
    instructions[4868] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149, 'op': 'addl'}
    instructions[4869] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149, 'op': 'addl'}
    instructions[4870] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149, 'op': 'addl'}
    instructions[4871] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149, 'op': 'load'}
    instructions[4872] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149, 'op': 'store'}
    instructions[4873] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149, 'op': 'addl'}
    instructions[4874] = {5'd0, 4'd8, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149 {'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149, 'op': 'literal'}
    instructions[4875] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4876] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149, 'op': 'load'}
    instructions[4877] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149, 'op': 'add'}
    instructions[4878] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149, 'op': 'addl'}
    instructions[4879] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149, 'op': 'load'}
    instructions[4880] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4881] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149, 'op': 'load'}
    instructions[4882] = {5'd13, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149, 'op': 'not_equal'}
    instructions[4883] = {5'd8, 4'd0, 4'd8, 16'd4902};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149 {'a': 8, 'label': 4902, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149, 'op': 'jmp_if_false'}
    instructions[4884] = {5'd0, 4'd8, 4'd0, 16'd65535};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149 {'literal': 65535, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149, 'op': 'literal'}
    instructions[4885] = {5'd3, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149 {'a': 8, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149, 'op': 'literal_hi'}
    instructions[4886] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149, 'op': 'store'}
    instructions[4887] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149, 'op': 'addl'}
    instructions[4888] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149, 'op': 'addl'}
    instructions[4889] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149, 'op': 'addl'}
    instructions[4890] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149, 'op': 'load'}
    instructions[4891] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149, 'op': 'store'}
    instructions[4892] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149, 'op': 'addl'}
    instructions[4893] = {5'd0, 4'd8, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149 {'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149, 'op': 'literal'}
    instructions[4894] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4895] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149, 'op': 'load'}
    instructions[4896] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149, 'op': 'add'}
    instructions[4897] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149, 'op': 'addl'}
    instructions[4898] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149, 'op': 'load'}
    instructions[4899] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4900] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149, 'op': 'load'}
    instructions[4901] = {5'd13, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149, 'op': 'not_equal'}
    instructions[4902] = {5'd8, 4'd0, 4'd8, 16'd4910};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149 {'a': 8, 'label': 4910, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149, 'op': 'jmp_if_false'}
    instructions[4903] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149, 'op': 'literal'}
    instructions[4904] = {5'd0, 4'd2, 4'd0, 16'd591};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149 {'literal': 591, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149, 'op': 'literal'}
    instructions[4905] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149, 'op': 'store'}
    instructions[4906] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149, 'op': 'addl'}
    instructions[4907] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149, 'op': 'addl'}
    instructions[4908] = {5'd16, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149, 'op': 'return'}
    instructions[4909] = {5'd10, 4'd0, 4'd0, 16'd4910};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149 {'label': 4910, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 149, 'op': 'goto'}
    instructions[4910] = {5'd0, 4'd8, 4'd0, 16'd2054};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 152 {'literal': 2054, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 152, 'op': 'literal'}
    instructions[4911] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 152 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 152, 'op': 'store'}
    instructions[4912] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 152 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 152, 'op': 'addl'}
    instructions[4913] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 152 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 152, 'op': 'addl'}
    instructions[4914] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 152 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 152, 'op': 'addl'}
    instructions[4915] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 152 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 152, 'op': 'load'}
    instructions[4916] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 152 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 152, 'op': 'store'}
    instructions[4917] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 152 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 152, 'op': 'addl'}
    instructions[4918] = {5'd0, 4'd8, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 152 {'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 152, 'op': 'literal'}
    instructions[4919] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 152 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 152, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4920] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 152 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 152, 'op': 'load'}
    instructions[4921] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 152 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 152, 'op': 'add'}
    instructions[4922] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 152 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 152, 'op': 'addl'}
    instructions[4923] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 152 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 152, 'op': 'load'}
    instructions[4924] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 152 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 152, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4925] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 152 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 152, 'op': 'load'}
    instructions[4926] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 152 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 152, 'op': 'equal'}
    instructions[4927] = {5'd8, 4'd0, 4'd8, 16'd5278};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 152 {'a': 8, 'label': 5278, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 152, 'op': 'jmp_if_false'}
    instructions[4928] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 154 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 154, 'op': 'literal'}
    instructions[4929] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 154 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 154, 'op': 'store'}
    instructions[4930] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 154 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 154, 'op': 'addl'}
    instructions[4931] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 154 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 154, 'op': 'addl'}
    instructions[4932] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 154 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 154, 'op': 'addl'}
    instructions[4933] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 154 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 154, 'op': 'load'}
    instructions[4934] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 154 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 154, 'op': 'store'}
    instructions[4935] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 154 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 154, 'op': 'addl'}
    instructions[4936] = {5'd0, 4'd8, 4'd0, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 154 {'literal': 10, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 154, 'op': 'literal'}
    instructions[4937] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 154 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 154, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4938] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 154 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 154, 'op': 'load'}
    instructions[4939] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 154 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 154, 'op': 'add'}
    instructions[4940] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 154 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 154, 'op': 'addl'}
    instructions[4941] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 154 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 154, 'op': 'load'}
    instructions[4942] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 154 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 154, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4943] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 154 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 154, 'op': 'load'}
    instructions[4944] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 154 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 154, 'op': 'equal'}
    instructions[4945] = {5'd8, 4'd0, 4'd8, 16'd5271};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 154 {'a': 8, 'label': 5271, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 154, 'op': 'jmp_if_false'}
    instructions[4946] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155, 'op': 'store'}
    instructions[4947] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155, 'op': 'addl'}
    instructions[4948] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155, 'op': 'store'}
    instructions[4949] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155, 'op': 'addl'}
    instructions[4950] = {5'd0, 4'd8, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155 {'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155, 'op': 'literal'}
    instructions[4951] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155, 'op': 'store'}
    instructions[4952] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155, 'op': 'addl'}
    instructions[4953] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155, 'op': 'addl'}
    instructions[4954] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155, 'op': 'addl'}
    instructions[4955] = {5'd4, 4'd6, 4'd0, 16'd5296};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155 {'z': 6, 'label': 5296, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155, 'op': 'call'}
    instructions[4956] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155, 'op': 'addl'}
    instructions[4957] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4958] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155, 'op': 'load'}
    instructions[4959] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4960] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155, 'op': 'load'}
    instructions[4961] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 155, 'op': 'addl'}
    instructions[4962] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 157 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 157, 'op': 'literal'}
    instructions[4963] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 157 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 157, 'op': 'store'}
    instructions[4964] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 157 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 157, 'op': 'addl'}
    instructions[4965] = {5'd0, 4'd8, 4'd0, 16'd27};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 157 {'literal': 27, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 157, 'op': 'literal'}
    instructions[4966] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 157 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 157, 'op': 'store'}
    instructions[4967] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 157 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 157, 'op': 'addl'}
    instructions[4968] = {5'd0, 4'd8, 4'd0, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 157 {'literal': 7, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 157, 'op': 'literal'}
    instructions[4969] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 157 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 157, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4970] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 157 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 157, 'op': 'load'}
    instructions[4971] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 157 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 157, 'op': 'add'}
    instructions[4972] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 157 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 157, 'op': 'addl'}
    instructions[4973] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 157 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 157, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4974] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 157 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 157, 'op': 'load'}
    instructions[4975] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 157 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 157, 'op': 'store'}
    instructions[4976] = {5'd0, 4'd8, 4'd0, 16'd2048};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 158 {'literal': 2048, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 158, 'op': 'literal'}
    instructions[4977] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 158 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 158, 'op': 'store'}
    instructions[4978] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 158 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 158, 'op': 'addl'}
    instructions[4979] = {5'd0, 4'd8, 4'd0, 16'd27};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 158 {'literal': 27, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 158, 'op': 'literal'}
    instructions[4980] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 158 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 158, 'op': 'store'}
    instructions[4981] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 158 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 158, 'op': 'addl'}
    instructions[4982] = {5'd0, 4'd8, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 158 {'literal': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 158, 'op': 'literal'}
    instructions[4983] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 158 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 158, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4984] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 158 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 158, 'op': 'load'}
    instructions[4985] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 158 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 158, 'op': 'add'}
    instructions[4986] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 158 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 158, 'op': 'addl'}
    instructions[4987] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 158 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 158, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4988] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 158 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 158, 'op': 'load'}
    instructions[4989] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 158 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 158, 'op': 'store'}
    instructions[4990] = {5'd0, 4'd8, 4'd0, 16'd1540};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 159 {'literal': 1540, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 159, 'op': 'literal'}
    instructions[4991] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 159 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 159, 'op': 'store'}
    instructions[4992] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 159 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 159, 'op': 'addl'}
    instructions[4993] = {5'd0, 4'd8, 4'd0, 16'd27};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 159 {'literal': 27, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 159, 'op': 'literal'}
    instructions[4994] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 159 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 159, 'op': 'store'}
    instructions[4995] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 159 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 159, 'op': 'addl'}
    instructions[4996] = {5'd0, 4'd8, 4'd0, 16'd9};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 159 {'literal': 9, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 159, 'op': 'literal'}
    instructions[4997] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 159 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 159, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4998] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 159 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 159, 'op': 'load'}
    instructions[4999] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 159 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 159, 'op': 'add'}
    instructions[5000] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 159 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 159, 'op': 'addl'}
    instructions[5001] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 159 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 159, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5002] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 159 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 159, 'op': 'load'}
    instructions[5003] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 159 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 159, 'op': 'store'}
    instructions[5004] = {5'd0, 4'd8, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 160 {'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 160, 'op': 'literal'}
    instructions[5005] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 160 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 160, 'op': 'store'}
    instructions[5006] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 160 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 160, 'op': 'addl'}
    instructions[5007] = {5'd0, 4'd8, 4'd0, 16'd27};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 160 {'literal': 27, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 160, 'op': 'literal'}
    instructions[5008] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 160 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 160, 'op': 'store'}
    instructions[5009] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 160 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 160, 'op': 'addl'}
    instructions[5010] = {5'd0, 4'd8, 4'd0, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 160 {'literal': 10, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 160, 'op': 'literal'}
    instructions[5011] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 160 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 160, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5012] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 160 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 160, 'op': 'load'}
    instructions[5013] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 160 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 160, 'op': 'add'}
    instructions[5014] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 160 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 160, 'op': 'addl'}
    instructions[5015] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 160 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 160, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5016] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 160 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 160, 'op': 'load'}
    instructions[5017] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 160 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 160, 'op': 'store'}
    instructions[5018] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 161 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 161, 'op': 'literal'}
    instructions[5019] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 161 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 161, 'op': 'store'}
    instructions[5020] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 161 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 161, 'op': 'addl'}
    instructions[5021] = {5'd0, 4'd8, 4'd0, 16'd27};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 161 {'literal': 27, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 161, 'op': 'literal'}
    instructions[5022] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 161 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 161, 'op': 'store'}
    instructions[5023] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 161 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 161, 'op': 'addl'}
    instructions[5024] = {5'd0, 4'd8, 4'd0, 16'd11};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 161 {'literal': 11, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 161, 'op': 'literal'}
    instructions[5025] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 161 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 161, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5026] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 161 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 161, 'op': 'load'}
    instructions[5027] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 161 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 161, 'op': 'add'}
    instructions[5028] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 161 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 161, 'op': 'addl'}
    instructions[5029] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 161 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 161, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5030] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 161 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 161, 'op': 'load'}
    instructions[5031] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 161 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 161, 'op': 'store'}
    instructions[5032] = {5'd0, 4'd8, 4'd0, 16'd515};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 162 {'literal': 515, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 162, 'op': 'literal'}
    instructions[5033] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 162 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 162, 'op': 'store'}
    instructions[5034] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 162 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 162, 'op': 'addl'}
    instructions[5035] = {5'd0, 4'd8, 4'd0, 16'd27};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 162 {'literal': 27, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 162, 'op': 'literal'}
    instructions[5036] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 162 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 162, 'op': 'store'}
    instructions[5037] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 162 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 162, 'op': 'addl'}
    instructions[5038] = {5'd0, 4'd8, 4'd0, 16'd12};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 162 {'literal': 12, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 162, 'op': 'literal'}
    instructions[5039] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 162 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 162, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5040] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 162 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 162, 'op': 'load'}
    instructions[5041] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 162 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 162, 'op': 'add'}
    instructions[5042] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 162 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 162, 'op': 'addl'}
    instructions[5043] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 162 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 162, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5044] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 162 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 162, 'op': 'load'}
    instructions[5045] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 162 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 162, 'op': 'store'}
    instructions[5046] = {5'd0, 4'd8, 4'd0, 16'd1029};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 163 {'literal': 1029, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 163, 'op': 'literal'}
    instructions[5047] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 163 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 163, 'op': 'store'}
    instructions[5048] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 163 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 163, 'op': 'addl'}
    instructions[5049] = {5'd0, 4'd8, 4'd0, 16'd27};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 163 {'literal': 27, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 163, 'op': 'literal'}
    instructions[5050] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 163 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 163, 'op': 'store'}
    instructions[5051] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 163 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 163, 'op': 'addl'}
    instructions[5052] = {5'd0, 4'd8, 4'd0, 16'd13};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 163 {'literal': 13, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 163, 'op': 'literal'}
    instructions[5053] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 163 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 163, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5054] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 163 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 163, 'op': 'load'}
    instructions[5055] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 163 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 163, 'op': 'add'}
    instructions[5056] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 163 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 163, 'op': 'addl'}
    instructions[5057] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 163 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 163, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5058] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 163 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 163, 'op': 'load'}
    instructions[5059] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 163 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 163, 'op': 'store'}
    instructions[5060] = {5'd0, 4'd8, 4'd0, 16'd49320};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 164 {'literal': 49320, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 164, 'op': 'literal'}
    instructions[5061] = {5'd3, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 164 {'a': 8, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 164, 'op': 'literal_hi'}
    instructions[5062] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 164 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 164, 'op': 'store'}
    instructions[5063] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 164 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 164, 'op': 'addl'}
    instructions[5064] = {5'd0, 4'd8, 4'd0, 16'd27};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 164 {'literal': 27, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 164, 'op': 'literal'}
    instructions[5065] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 164 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 164, 'op': 'store'}
    instructions[5066] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 164 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 164, 'op': 'addl'}
    instructions[5067] = {5'd0, 4'd8, 4'd0, 16'd14};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 164 {'literal': 14, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 164, 'op': 'literal'}
    instructions[5068] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 164 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 164, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5069] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 164 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 164, 'op': 'load'}
    instructions[5070] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 164 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 164, 'op': 'add'}
    instructions[5071] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 164 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 164, 'op': 'addl'}
    instructions[5072] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 164 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 164, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5073] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 164 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 164, 'op': 'load'}
    instructions[5074] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 164 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 164, 'op': 'store'}
    instructions[5075] = {5'd0, 4'd8, 4'd0, 16'd257};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 165 {'literal': 257, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 165, 'op': 'literal'}
    instructions[5076] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 165 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 165, 'op': 'store'}
    instructions[5077] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 165 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 165, 'op': 'addl'}
    instructions[5078] = {5'd0, 4'd8, 4'd0, 16'd27};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 165 {'literal': 27, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 165, 'op': 'literal'}
    instructions[5079] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 165 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 165, 'op': 'store'}
    instructions[5080] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 165 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 165, 'op': 'addl'}
    instructions[5081] = {5'd0, 4'd8, 4'd0, 16'd15};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 165 {'literal': 15, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 165, 'op': 'literal'}
    instructions[5082] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 165 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 165, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5083] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 165 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 165, 'op': 'load'}
    instructions[5084] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 165 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 165, 'op': 'add'}
    instructions[5085] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 165 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 165, 'op': 'addl'}
    instructions[5086] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 165 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 165, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5087] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 165 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 165, 'op': 'load'}
    instructions[5088] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 165 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 165, 'op': 'store'}
    instructions[5089] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166, 'op': 'addl'}
    instructions[5090] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166, 'op': 'addl'}
    instructions[5091] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166, 'op': 'load'}
    instructions[5092] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166, 'op': 'store'}
    instructions[5093] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166, 'op': 'addl'}
    instructions[5094] = {5'd0, 4'd8, 4'd0, 16'd11};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166 {'literal': 11, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166, 'op': 'literal'}
    instructions[5095] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5096] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166, 'op': 'load'}
    instructions[5097] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166, 'op': 'add'}
    instructions[5098] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166, 'op': 'addl'}
    instructions[5099] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166, 'op': 'load'}
    instructions[5100] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166, 'op': 'store'}
    instructions[5101] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166, 'op': 'addl'}
    instructions[5102] = {5'd0, 4'd8, 4'd0, 16'd27};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166 {'literal': 27, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166, 'op': 'literal'}
    instructions[5103] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166, 'op': 'store'}
    instructions[5104] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166, 'op': 'addl'}
    instructions[5105] = {5'd0, 4'd8, 4'd0, 16'd16};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166 {'literal': 16, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166, 'op': 'literal'}
    instructions[5106] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5107] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166, 'op': 'load'}
    instructions[5108] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166, 'op': 'add'}
    instructions[5109] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166, 'op': 'addl'}
    instructions[5110] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5111] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166, 'op': 'load'}
    instructions[5112] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 166, 'op': 'store'}
    instructions[5113] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167, 'op': 'addl'}
    instructions[5114] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167, 'op': 'addl'}
    instructions[5115] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167, 'op': 'load'}
    instructions[5116] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167, 'op': 'store'}
    instructions[5117] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167, 'op': 'addl'}
    instructions[5118] = {5'd0, 4'd8, 4'd0, 16'd12};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167 {'literal': 12, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167, 'op': 'literal'}
    instructions[5119] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5120] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167, 'op': 'load'}
    instructions[5121] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167, 'op': 'add'}
    instructions[5122] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167, 'op': 'addl'}
    instructions[5123] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167, 'op': 'load'}
    instructions[5124] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167, 'op': 'store'}
    instructions[5125] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167, 'op': 'addl'}
    instructions[5126] = {5'd0, 4'd8, 4'd0, 16'd27};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167 {'literal': 27, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167, 'op': 'literal'}
    instructions[5127] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167, 'op': 'store'}
    instructions[5128] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167, 'op': 'addl'}
    instructions[5129] = {5'd0, 4'd8, 4'd0, 16'd17};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167 {'literal': 17, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167, 'op': 'literal'}
    instructions[5130] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5131] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167, 'op': 'load'}
    instructions[5132] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167, 'op': 'add'}
    instructions[5133] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167, 'op': 'addl'}
    instructions[5134] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5135] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167, 'op': 'load'}
    instructions[5136] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 167, 'op': 'store'}
    instructions[5137] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168, 'op': 'addl'}
    instructions[5138] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168, 'op': 'addl'}
    instructions[5139] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168, 'op': 'load'}
    instructions[5140] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168, 'op': 'store'}
    instructions[5141] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168, 'op': 'addl'}
    instructions[5142] = {5'd0, 4'd8, 4'd0, 16'd13};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168 {'literal': 13, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168, 'op': 'literal'}
    instructions[5143] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5144] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168, 'op': 'load'}
    instructions[5145] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168, 'op': 'add'}
    instructions[5146] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168, 'op': 'addl'}
    instructions[5147] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168, 'op': 'load'}
    instructions[5148] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168, 'op': 'store'}
    instructions[5149] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168, 'op': 'addl'}
    instructions[5150] = {5'd0, 4'd8, 4'd0, 16'd27};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168 {'literal': 27, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168, 'op': 'literal'}
    instructions[5151] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168, 'op': 'store'}
    instructions[5152] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168, 'op': 'addl'}
    instructions[5153] = {5'd0, 4'd8, 4'd0, 16'd18};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168 {'literal': 18, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168, 'op': 'literal'}
    instructions[5154] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5155] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168, 'op': 'load'}
    instructions[5156] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168, 'op': 'add'}
    instructions[5157] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168, 'op': 'addl'}
    instructions[5158] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5159] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168, 'op': 'load'}
    instructions[5160] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 168, 'op': 'store'}
    instructions[5161] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169, 'op': 'addl'}
    instructions[5162] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169, 'op': 'addl'}
    instructions[5163] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169, 'op': 'load'}
    instructions[5164] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169, 'op': 'store'}
    instructions[5165] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169, 'op': 'addl'}
    instructions[5166] = {5'd0, 4'd8, 4'd0, 16'd14};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169 {'literal': 14, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169, 'op': 'literal'}
    instructions[5167] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5168] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169, 'op': 'load'}
    instructions[5169] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169, 'op': 'add'}
    instructions[5170] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169, 'op': 'addl'}
    instructions[5171] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169, 'op': 'load'}
    instructions[5172] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169, 'op': 'store'}
    instructions[5173] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169, 'op': 'addl'}
    instructions[5174] = {5'd0, 4'd8, 4'd0, 16'd27};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169 {'literal': 27, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169, 'op': 'literal'}
    instructions[5175] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169, 'op': 'store'}
    instructions[5176] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169, 'op': 'addl'}
    instructions[5177] = {5'd0, 4'd8, 4'd0, 16'd19};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169 {'literal': 19, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169, 'op': 'literal'}
    instructions[5178] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5179] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169, 'op': 'load'}
    instructions[5180] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169, 'op': 'add'}
    instructions[5181] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169, 'op': 'addl'}
    instructions[5182] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5183] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169, 'op': 'load'}
    instructions[5184] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 169, 'op': 'store'}
    instructions[5185] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170, 'op': 'addl'}
    instructions[5186] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170, 'op': 'addl'}
    instructions[5187] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170, 'op': 'load'}
    instructions[5188] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170, 'op': 'store'}
    instructions[5189] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170, 'op': 'addl'}
    instructions[5190] = {5'd0, 4'd8, 4'd0, 16'd15};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170 {'literal': 15, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170, 'op': 'literal'}
    instructions[5191] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5192] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170, 'op': 'load'}
    instructions[5193] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170, 'op': 'add'}
    instructions[5194] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170, 'op': 'addl'}
    instructions[5195] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170, 'op': 'load'}
    instructions[5196] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170, 'op': 'store'}
    instructions[5197] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170, 'op': 'addl'}
    instructions[5198] = {5'd0, 4'd8, 4'd0, 16'd27};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170 {'literal': 27, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170, 'op': 'literal'}
    instructions[5199] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170, 'op': 'store'}
    instructions[5200] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170, 'op': 'addl'}
    instructions[5201] = {5'd0, 4'd8, 4'd0, 16'd20};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170 {'literal': 20, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170, 'op': 'literal'}
    instructions[5202] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5203] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170, 'op': 'load'}
    instructions[5204] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170, 'op': 'add'}
    instructions[5205] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170, 'op': 'addl'}
    instructions[5206] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5207] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170, 'op': 'load'}
    instructions[5208] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 170, 'op': 'store'}
    instructions[5209] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171, 'op': 'store'}
    instructions[5210] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171, 'op': 'addl'}
    instructions[5211] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171, 'op': 'store'}
    instructions[5212] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171, 'op': 'addl'}
    instructions[5213] = {5'd0, 4'd8, 4'd0, 16'd27};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 172 {'literal': 27, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 172, 'op': 'literal'}
    instructions[5214] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171, 'op': 'store'}
    instructions[5215] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171, 'op': 'addl'}
    instructions[5216] = {5'd0, 4'd8, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 173 {'literal': 60, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 173, 'op': 'literal'}
    instructions[5217] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171, 'op': 'store'}
    instructions[5218] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171, 'op': 'addl'}
    instructions[5219] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 174 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 174, 'op': 'addl'}
    instructions[5220] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 174 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 174, 'op': 'addl'}
    instructions[5221] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 174 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 174, 'op': 'load'}
    instructions[5222] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 174 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 174, 'op': 'store'}
    instructions[5223] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 174 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 174, 'op': 'addl'}
    instructions[5224] = {5'd0, 4'd8, 4'd0, 16'd11};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 174 {'literal': 11, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 174, 'op': 'literal'}
    instructions[5225] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 174 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 174, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5226] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 174 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 174, 'op': 'load'}
    instructions[5227] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 174 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 174, 'op': 'add'}
    instructions[5228] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 174 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 174, 'op': 'addl'}
    instructions[5229] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 174 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 174, 'op': 'load'}
    instructions[5230] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171, 'op': 'store'}
    instructions[5231] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171, 'op': 'addl'}
    instructions[5232] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 175 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 175, 'op': 'addl'}
    instructions[5233] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 175 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 175, 'op': 'addl'}
    instructions[5234] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 175 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 175, 'op': 'load'}
    instructions[5235] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 175 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 175, 'op': 'store'}
    instructions[5236] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 175 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 175, 'op': 'addl'}
    instructions[5237] = {5'd0, 4'd8, 4'd0, 16'd12};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 175 {'literal': 12, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 175, 'op': 'literal'}
    instructions[5238] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 175 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 175, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5239] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 175 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 175, 'op': 'load'}
    instructions[5240] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 175 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 175, 'op': 'add'}
    instructions[5241] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 175 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 175, 'op': 'addl'}
    instructions[5242] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 175 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 175, 'op': 'load'}
    instructions[5243] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171, 'op': 'store'}
    instructions[5244] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171, 'op': 'addl'}
    instructions[5245] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 176 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 176, 'op': 'addl'}
    instructions[5246] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 176 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 176, 'op': 'addl'}
    instructions[5247] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 176 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 176, 'op': 'load'}
    instructions[5248] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 176 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 176, 'op': 'store'}
    instructions[5249] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 176 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 176, 'op': 'addl'}
    instructions[5250] = {5'd0, 4'd8, 4'd0, 16'd13};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 176 {'literal': 13, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 176, 'op': 'literal'}
    instructions[5251] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 176 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 176, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5252] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 176 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 176, 'op': 'load'}
    instructions[5253] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 176 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 176, 'op': 'add'}
    instructions[5254] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 176 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 176, 'op': 'addl'}
    instructions[5255] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 176 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 176, 'op': 'load'}
    instructions[5256] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171, 'op': 'store'}
    instructions[5257] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171, 'op': 'addl'}
    instructions[5258] = {5'd0, 4'd8, 4'd0, 16'd2054};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 177 {'literal': 2054, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 177, 'op': 'literal'}
    instructions[5259] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171, 'op': 'store'}
    instructions[5260] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171, 'op': 'addl'}
    instructions[5261] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171, 'op': 'addl'}
    instructions[5262] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171, 'op': 'addl'}
    instructions[5263] = {5'd4, 4'd6, 4'd0, 16'd3081};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171 {'z': 6, 'label': 3081, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171, 'op': 'call'}
    instructions[5264] = {5'd1, 4'd3, 4'd3, -16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171 {'a': 3, 'literal': -6, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171, 'op': 'addl'}
    instructions[5265] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5266] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171, 'op': 'load'}
    instructions[5267] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5268] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171, 'op': 'load'}
    instructions[5269] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 171, 'op': 'addl'}
    instructions[5270] = {5'd10, 4'd0, 4'd0, 16'd5271};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 154 {'label': 5271, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 154, 'op': 'goto'}
    instructions[5271] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 179 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 179, 'op': 'literal'}
    instructions[5272] = {5'd0, 4'd2, 4'd0, 16'd591};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 179 {'literal': 591, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 179, 'op': 'literal'}
    instructions[5273] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 179 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 179, 'op': 'store'}
    instructions[5274] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 179 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 179, 'op': 'addl'}
    instructions[5275] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 179 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 179, 'op': 'addl'}
    instructions[5276] = {5'd16, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 179 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 179, 'op': 'return'}
    instructions[5277] = {5'd10, 4'd0, 4'd0, 16'd5278};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 152 {'label': 5278, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 152, 'op': 'goto'}
    instructions[5278] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 181 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 181, 'op': 'addl'}
    instructions[5279] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 181 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 181, 'op': 'addl'}
    instructions[5280] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 181 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 181, 'op': 'load'}
    instructions[5281] = {5'd0, 4'd2, 4'd0, 16'd591};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 181 {'literal': 591, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 181, 'op': 'literal'}
    instructions[5282] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 181 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 181, 'op': 'store'}
    instructions[5283] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 181 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 181, 'op': 'addl'}
    instructions[5284] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 181 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 181, 'op': 'addl'}
    instructions[5285] = {5'd16, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 181 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 181, 'op': 'return'}
    instructions[5286] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 27 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 27, 'op': 'addl'}
    instructions[5287] = {5'd0, 4'd8, 4'd0, 16'd654};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 28 {'literal': 654, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 28, 'op': 'literal'}
    instructions[5288] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 28 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 28, 'op': 'addl'}
    instructions[5289] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 28 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 28, 'op': 'load'}
    instructions[5290] = {5'd14, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 28 {'a': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 28, 'op': 'ready'}
    instructions[5291] = {5'd0, 4'd2, 4'd0, 16'd26};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 28 {'literal': 26, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 28, 'op': 'literal'}
    instructions[5292] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 28 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 28, 'op': 'store'}
    instructions[5293] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 28 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 28, 'op': 'addl'}
    instructions[5294] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 28 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 28, 'op': 'addl'}
    instructions[5295] = {5'd16, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 28 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 28, 'op': 'return'}
    instructions[5296] = {5'd1, 4'd3, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73 {'a': 3, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73, 'op': 'addl'}
    instructions[5297] = {5'd2, 4'd0, 4'd3, 16'd6};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'store'}
    instructions[5298] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[5299] = {5'd2, 4'd0, 4'd3, 16'd7};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'store'}
    instructions[5300] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[5301] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[5302] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[5303] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'load'}
    instructions[5304] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'store'}
    instructions[5305] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[5306] = {5'd0, 4'd8, 4'd0, 16'd24};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'literal': 24, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'literal'}
    instructions[5307] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[5308] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'load'}
    instructions[5309] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'store'}
    instructions[5310] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[5311] = {5'd1, 4'd7, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 4, 'literal': 0, 'z': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[5312] = {5'd1, 4'd4, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[5313] = {5'd4, 4'd6, 4'd0, 16'd5323};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'z': 6, 'label': 5323, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'call'}
    instructions[5314] = {5'd1, 4'd3, 4'd3, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': -2, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[5315] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5316] = {5'd6, 4'd7, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'z': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'load'}
    instructions[5317] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5318] = {5'd6, 4'd6, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'z': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'load'}
    instructions[5319] = {5'd1, 4'd3, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[5320] = {5'd1, 4'd3, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73 {'a': 4, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73, 'op': 'addl'}
    instructions[5321] = {5'd1, 4'd4, 4'd7, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73 {'a': 7, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73, 'op': 'addl'}
    instructions[5322] = {5'd16, 4'd0, 4'd6, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73 {'a': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73, 'op': 'return'}
    instructions[5323] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23, 'op': 'addl'}
    instructions[5324] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 24 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 24, 'op': 'literal'}
    instructions[5325] = {5'd1, 4'd2, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 24 {'a': 4, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 24, 'op': 'addl'}
    instructions[5326] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 24 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 24, 'op': 'store'}
    instructions[5327] = {5'd1, 4'd8, 4'd4, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 4, 'literal': -2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'addl'}
    instructions[5328] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'addl'}
    instructions[5329] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'load'}
    instructions[5330] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'store'}
    instructions[5331] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'addl'}
    instructions[5332] = {5'd1, 4'd8, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 4, 'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'addl'}
    instructions[5333] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'addl'}
    instructions[5334] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'load'}
    instructions[5335] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5336] = {5'd6, 4'd2, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 3, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'load'}
    instructions[5337] = {5'd7, 4'd8, 4'd8, 16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 8, 'z': 8, 'b': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'add'}
    instructions[5338] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'addl'}
    instructions[5339] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'load'}
    instructions[5340] = {5'd8, 4'd0, 4'd8, 16'd5382};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 29 {'a': 8, 'label': 5382, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 29, 'op': 'jmp_if_false'}
    instructions[5341] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[5342] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[5343] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'load'}
    instructions[5344] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'store'}
    instructions[5345] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[5346] = {5'd1, 4'd8, 4'd4, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 4, 'literal': -2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[5347] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[5348] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'load'}
    instructions[5349] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'store'}
    instructions[5350] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[5351] = {5'd1, 4'd8, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 4, 'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[5352] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[5353] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'load'}
    instructions[5354] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5355] = {5'd6, 4'd2, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'load'}
    instructions[5356] = {5'd7, 4'd8, 4'd8, 16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 8, 'z': 8, 'b': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'add'}
    instructions[5357] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[5358] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'load'}
    instructions[5359] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5360] = {5'd6, 4'd0, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'z': 0, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'load'}
    instructions[5361] = {5'd25, 4'd0, 4'd0, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 0, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'write'}
    instructions[5362] = {5'd1, 4'd3, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[5363] = {5'd1, 4'd8, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 4, 'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[5364] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[5365] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'load'}
    instructions[5366] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'store'}
    instructions[5367] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[5368] = {5'd0, 4'd8, 4'd0, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'literal': 1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'literal'}
    instructions[5369] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'store'}
    instructions[5370] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[5371] = {5'd1, 4'd8, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 4, 'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[5372] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[5373] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'load'}
    instructions[5374] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5375] = {5'd6, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'load'}
    instructions[5376] = {5'd7, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'add'}
    instructions[5377] = {5'd1, 4'd2, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 4, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[5378] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'store'}
    instructions[5379] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5380] = {5'd6, 4'd8, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'load'}
    instructions[5381] = {5'd10, 4'd0, 4'd0, 16'd5383};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 29 {'label': 5383, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 29, 'op': 'goto'}
    instructions[5382] = {5'd10, 4'd0, 4'd0, 16'd5384};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 29 {'label': 5384, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 29, 'op': 'goto'}
    instructions[5383] = {5'd10, 4'd0, 4'd0, 16'd5327};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'label': 5327, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'goto'}
    instructions[5384] = {5'd1, 4'd3, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23 {'a': 4, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23, 'op': 'addl'}
    instructions[5385] = {5'd1, 4'd4, 4'd7, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23 {'a': 7, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23, 'op': 'addl'}
    instructions[5386] = {5'd16, 4'd0, 4'd6, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23 {'a': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23, 'op': 'return'}
    instructions[5387] = {5'd1, 4'd3, 4'd3, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 481 {'a': 3, 'literal': 2, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 481, 'op': 'addl'}
    instructions[5388] = {5'd1, 4'd8, 4'd4, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 484 {'a': 4, 'literal': -2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 484, 'op': 'addl'}
    instructions[5389] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 484 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 484, 'op': 'addl'}
    instructions[5390] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 484 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 484, 'op': 'load'}
    instructions[5391] = {5'd1, 4'd2, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 484 {'a': 4, 'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 484, 'op': 'addl'}
    instructions[5392] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 484 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 484, 'op': 'store'}
    instructions[5393] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 485 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 485, 'op': 'store'}
    instructions[5394] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 485 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 485, 'op': 'addl'}
    instructions[5395] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 485 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 485, 'op': 'store'}
    instructions[5396] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 485 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 485, 'op': 'addl'}
    instructions[5397] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 485 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 485, 'op': 'addl'}
    instructions[5398] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 485 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 485, 'op': 'addl'}
    instructions[5399] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 485 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 485, 'op': 'load'}
    instructions[5400] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 485 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 485, 'op': 'store'}
    instructions[5401] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 485 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 485, 'op': 'addl'}
    instructions[5402] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 485 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 485, 'op': 'addl'}
    instructions[5403] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 485 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 485, 'op': 'addl'}
    instructions[5404] = {5'd4, 4'd6, 4'd0, 16'd5487};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 485 {'z': 6, 'label': 5487, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 485, 'op': 'call'}
    instructions[5405] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 485 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 485, 'op': 'addl'}
    instructions[5406] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 485 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 485, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5407] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 485 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 485, 'op': 'load'}
    instructions[5408] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 485 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 485, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5409] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 485 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 485, 'op': 'load'}
    instructions[5410] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 485 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 485, 'op': 'addl'}
    instructions[5411] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486, 'op': 'literal'}
    instructions[5412] = {5'd1, 4'd2, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486, 'op': 'addl'}
    instructions[5413] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486, 'op': 'store'}
    instructions[5414] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486, 'op': 'addl'}
    instructions[5415] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486, 'op': 'addl'}
    instructions[5416] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486, 'op': 'load'}
    instructions[5417] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486, 'op': 'store'}
    instructions[5418] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486, 'op': 'addl'}
    instructions[5419] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486, 'op': 'addl'}
    instructions[5420] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486, 'op': 'addl'}
    instructions[5421] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486, 'op': 'load'}
    instructions[5422] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5423] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486, 'op': 'load'}
    instructions[5424] = {5'd19, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486, 'op': 'unsigned_greater'}
    instructions[5425] = {5'd8, 4'd0, 4'd8, 16'd5484};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486 {'a': 8, 'label': 5484, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486, 'op': 'jmp_if_false'}
    instructions[5426] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487, 'op': 'store'}
    instructions[5427] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487, 'op': 'addl'}
    instructions[5428] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487, 'op': 'store'}
    instructions[5429] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487, 'op': 'addl'}
    instructions[5430] = {5'd1, 4'd8, 4'd4, -16'd3};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487 {'a': 4, 'literal': -3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487, 'op': 'addl'}
    instructions[5431] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487, 'op': 'addl'}
    instructions[5432] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487, 'op': 'load'}
    instructions[5433] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487, 'op': 'store'}
    instructions[5434] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487, 'op': 'addl'}
    instructions[5435] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487, 'op': 'addl'}
    instructions[5436] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487, 'op': 'addl'}
    instructions[5437] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487, 'op': 'load'}
    instructions[5438] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5439] = {5'd6, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487, 'op': 'load'}
    instructions[5440] = {5'd7, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487, 'op': 'add'}
    instructions[5441] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487, 'op': 'addl'}
    instructions[5442] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487, 'op': 'load'}
    instructions[5443] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487, 'op': 'store'}
    instructions[5444] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487, 'op': 'addl'}
    instructions[5445] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487, 'op': 'addl'}
    instructions[5446] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487, 'op': 'addl'}
    instructions[5447] = {5'd4, 4'd6, 4'd0, 16'd5487};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487 {'z': 6, 'label': 5487, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487, 'op': 'call'}
    instructions[5448] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487, 'op': 'addl'}
    instructions[5449] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5450] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487, 'op': 'load'}
    instructions[5451] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5452] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487, 'op': 'load'}
    instructions[5453] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 487, 'op': 'addl'}
    instructions[5454] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 488 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 488, 'op': 'addl'}
    instructions[5455] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 488 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 488, 'op': 'addl'}
    instructions[5456] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 488 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 488, 'op': 'load'}
    instructions[5457] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 488 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 488, 'op': 'store'}
    instructions[5458] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 488 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 488, 'op': 'addl'}
    instructions[5459] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 488 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 488, 'op': 'literal'}
    instructions[5460] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 488 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 488, 'op': 'store'}
    instructions[5461] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 488 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 488, 'op': 'addl'}
    instructions[5462] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 488 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 488, 'op': 'addl'}
    instructions[5463] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 488 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 488, 'op': 'addl'}
    instructions[5464] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 488 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 488, 'op': 'load'}
    instructions[5465] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 488 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 488, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5466] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 488 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 488, 'op': 'load'}
    instructions[5467] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 488 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 488, 'op': 'add'}
    instructions[5468] = {5'd1, 4'd2, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 488 {'a': 4, 'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 488, 'op': 'addl'}
    instructions[5469] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 488 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 488, 'op': 'store'}
    instructions[5470] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 488 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 488, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5471] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 488 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 488, 'op': 'load'}
    instructions[5472] = {5'd0, 4'd8, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486 {'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486, 'op': 'literal'}
    instructions[5473] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486, 'op': 'store'}
    instructions[5474] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486, 'op': 'addl'}
    instructions[5475] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486, 'op': 'addl'}
    instructions[5476] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486, 'op': 'addl'}
    instructions[5477] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486, 'op': 'load'}
    instructions[5478] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5479] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486, 'op': 'load'}
    instructions[5480] = {5'd7, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486, 'op': 'add'}
    instructions[5481] = {5'd1, 4'd2, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486, 'op': 'addl'}
    instructions[5482] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486, 'op': 'store'}
    instructions[5483] = {5'd10, 4'd0, 4'd0, 16'd5414};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486 {'label': 5414, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 486, 'op': 'goto'}
    instructions[5484] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 481 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 481, 'op': 'addl'}
    instructions[5485] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 481 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 481, 'op': 'addl'}
    instructions[5486] = {5'd16, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 481 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 481, 'op': 'return'}
    instructions[5487] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 21 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 21, 'op': 'addl'}
    instructions[5488] = {5'd0, 4'd8, 4'd0, 16'd544};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 22 {'literal': 544, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 22, 'op': 'literal'}
    instructions[5489] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 22 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 22, 'op': 'addl'}
    instructions[5490] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 22 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 22, 'op': 'load'}
    instructions[5491] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 22 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 22, 'op': 'store'}
    instructions[5492] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 22 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 22, 'op': 'addl'}
    instructions[5493] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 22 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 22, 'op': 'addl'}
    instructions[5494] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 22 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 22, 'op': 'addl'}
    instructions[5495] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 22 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 22, 'op': 'load'}
    instructions[5496] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 22 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 22, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5497] = {5'd6, 4'd0, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 22 {'a': 3, 'z': 0, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 22, 'op': 'load'}
    instructions[5498] = {5'd25, 4'd0, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 22 {'a': 0, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 22, 'op': 'write'}
    instructions[5499] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 22 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 22, 'op': 'addl'}
    instructions[5500] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 21 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 21, 'op': 'addl'}
    instructions[5501] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 21 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 21, 'op': 'addl'}
    instructions[5502] = {5'd16, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 21 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/web_server/server.c : 21, 'op': 'return'}
  end

  
  always @(posedge clk)
  begin
    load_data <= memory[load_address];
    if(store_enable && state == execute) begin
      memory[store_address] <= store_data;
    end
  end


  //////////////////////////////////////////////////////////////////////////////
  // PIPELINE STAGE 1 -- FETCH INSTRUCTION
  //                                                                            
  
  always @(posedge clk)
  begin
    //implement memory for instructions
    if (state == instruction_fetch || state == operand_fetch || state == execute) begin
      instruction <= instructions[program_counter];
      program_counter_1 <= program_counter;
    end
  end

  assign opcode    = instruction[28:24];
  assign address_z = instruction[23:20];
  assign address_a = instruction[19:16];
  assign address_b = instruction[3:0];
  assign literal   = instruction[15:0];

  //////////////////////////////////////////////////////////////////////////////
  // PIPELINE STAGE 2 -- FETCH OPERANDS
  //                                                                            
  
  always @(posedge clk)
  begin
    if (write_enable) begin
      registers[address_z_3] <= result;
    end
    if (state == operand_fetch || state == execute) begin
      opcode_2 <= opcode;
      literal_2 <= literal;
      address_a_2 <= address_a;
      address_b_2 <= address_b;
      address_z_2 <= address_z;
      program_counter_2 <= program_counter_1;
    end
  end
  assign register_a = registers[address_a_2];
  assign register_b = registers[address_b_2];
  assign operand_a = (address_a_2 == address_z_3 && write_enable)?result:register_a;
  assign operand_b = (address_b_2 == address_z_3 && write_enable)?result:register_b;
  assign store_address = operand_a;
  assign load_address = operand_a;
  assign store_data = operand_b;
  assign store_enable = (opcode_2==2);

  //////////////////////////////////////////////////////////////////////////////
  // PIPELINE STAGE 3 -- EXECUTE
  //                                                                            
  
  always @(posedge clk)
  begin

  write_enable <= 0;
  timer_clock <= timer_clock + 1;
  case(state)

    //instruction_fetch
    instruction_fetch: begin
      program_counter <= program_counter + 1;
      state <= operand_fetch;
    end
    //operand_fetch
    operand_fetch: begin
      program_counter <= program_counter + 1;
      state <= execute;
    end
    //execute
    execute: begin
      program_counter <= program_counter + 1;
      address_z_3 <= address_z_2;
      case(opcode_2)

        //literal
        16'd0:
        begin
          result<=$signed(literal_2);
          write_enable <= 1;
        end

        //addl
        16'd1:
        begin
          result<=operand_a + literal_2;
          write_enable <= 1;
        end

        //store
        16'd2:
        begin
        end

        //literal_hi
        16'd3:
        begin
          result<= {literal_2, operand_a[15:0]};
          write_enable <= 1;
        end

        //call
        16'd4:
        begin
          result <= program_counter_2 + 1;
          write_enable <= 1;
          program_counter <= literal_2;
          state <= instruction_fetch;
        end

        //stop
        16'd5:
        begin
        state <= stop;
        end

        //load
        16'd6:
        begin
          state <= load;
        end

        //add
        16'd7:
        begin
          long_result = operand_a + operand_b;
          result <= long_result[31:0];
          carry[0] <= long_result[32];
          write_enable <= 1;
        end

        //jmp_if_false
        16'd8:
        begin
          if (operand_a == 0) begin
            program_counter <= literal_2;
            state <= instruction_fetch;
          end
        end

        //subtract
        16'd9:
        begin
          long_result = operand_a + (~operand_b) + 1;
          result <= long_result[31:0];
          carry[0] <= ~long_result[32];
          write_enable <= 1;
        end

        //goto
        16'd10:
        begin
          program_counter <= literal_2;
          state <= instruction_fetch;
        end

        //equal
        16'd11:
        begin
          result <= operand_a == operand_b;
          write_enable <= 1;
        end

        //jmp_if_true
        16'd12:
        begin
          if (operand_a != 0) begin
            program_counter <= literal_2;
            state <= instruction_fetch;
          end
        end

        //not_equal
        16'd13:
        begin
          result <= operand_a != operand_b;
          write_enable <= 1;
        end

        //ready
        16'd14:
        begin
          result <= 0;
          case(operand_a)

            2:
            begin
              result[0] <= input_eth_rx_stb;
            end
            3:
            begin
              result[0] <= input_socket_stb;
            end
          endcase
          write_enable <= 1;
        end

        //wait_clocks
        16'd15:
        begin
          timer <= operand_a;
          state <= wait_state;
        end

        //return
        16'd16:
        begin
          program_counter <= operand_a;
          state <= instruction_fetch;
        end

        //or
        16'd17:
        begin
          result <= operand_a | operand_b;
          write_enable <= 1;
        end

        //unsigned_shift_right
        16'd18:
        begin
          if(operand_b < 32) begin
            result <= operand_a >> operand_b;
            carry <= operand_a << (32-operand_b);
          end else begin
            result <= 0;
            carry <= operand_a;
          end
          write_enable <= 1;
        end

        //unsigned_greater
        16'd19:
        begin
          result <= $unsigned(operand_a) > $unsigned(operand_b);
          write_enable <= 1;
        end

        //int_to_long
        16'd20:
        begin
          if(operand_a[31]) begin
            result <= -1;
          end else begin
            result <= 0;
          end
          write_enable <= 1;
        end

        //add_with_carry
        16'd21:
        begin
          long_result = operand_a + operand_b + carry[0];
          result <= long_result[31:0];
          carry[0] <= long_result[32];
          write_enable <= 1;
        end

        //and
        16'd22:
        begin
          result <= operand_a & operand_b;
          write_enable <= 1;
        end

        //not
        16'd23:
        begin
          result <= ~operand_a;
          write_enable <= 1;
        end

        //unsigned_greater_equal
        16'd24:
        begin
          result <= $unsigned(operand_a) >= $unsigned(operand_b);
          write_enable <= 1;
        end

        //write
        16'd25:
        begin
          state <= write;
          write_output <= operand_a;
          write_value <= operand_b;
        end

        //read
        16'd26:
        begin
          state <= read;
          read_input <= operand_a;
        end

        //shift_right
        16'd27:
        begin
          if(operand_b < 32) begin
            result <= $signed(operand_a) >>> operand_b;
            carry <= operand_a << (32-operand_b);
          end else begin
            result <= operand_a[31]?-1:0;
            carry <= operand_a;
          end
          write_enable <= 1;
        end

        //shift_left
        16'd28:
        begin
          if(operand_b < 32) begin
            result <= operand_a << operand_b;
            carry <= operand_a >> (32-operand_b);
          end else begin
            result <= 0;
            carry <= operand_a;
          end
          write_enable <= 1;
        end

      endcase

    end

    read:
    begin
      case(read_input)
      2:
      begin
        s_input_eth_rx_ack <= 1;
        if (s_input_eth_rx_ack && input_eth_rx_stb) begin
          result <= input_eth_rx;
          write_enable <= 1;
          s_input_eth_rx_ack <= 0;
          state <= execute;
        end
      end
      3:
      begin
        s_input_socket_ack <= 1;
        if (s_input_socket_ack && input_socket_stb) begin
          result <= input_socket;
          write_enable <= 1;
          s_input_socket_ack <= 0;
          state <= execute;
        end
      end
      endcase
    end

    write:
    begin
      case(write_output)
      0:
      begin
        s_output_eth_tx_stb <= 1;
        s_output_eth_tx <= write_value;
        if (output_eth_tx_ack && s_output_eth_tx_stb) begin
          s_output_eth_tx_stb <= 0;
          state <= execute;
        end
      end
      1:
      begin
        s_output_socket_stb <= 1;
        s_output_socket <= write_value;
        if (output_socket_ack && s_output_socket_stb) begin
          s_output_socket_stb <= 0;
          state <= execute;
        end
      end
      4:
      begin
        s_output_rs232_tx_stb <= 1;
        s_output_rs232_tx <= write_value;
        if (output_rs232_tx_ack && s_output_rs232_tx_stb) begin
          s_output_rs232_tx_stb <= 0;
          state <= execute;
        end
      end
      endcase
    end

    load:
    begin
        result <= load_data;
        write_enable <= 1;
        state <= execute;
    end

    wait_state:
    begin
      if (timer) begin
        timer <= timer - 1;
      end else begin
        state <= execute;
      end
    end

    stop:
    begin
    end

    endcase

    if (rst == 1'b1) begin
      timer <= 0;
      timer_clock <= 0;
      program_counter <= 0;
      address_z_3 <= 0;
      result <= 0;
      a = 0;
      b = 0;
      z = 0;
      state <= instruction_fetch;
      s_input_eth_rx_ack <= 0;
      s_input_socket_ack <= 0;
      s_output_eth_tx_stb <= 0;
      s_output_socket_stb <= 0;
      s_output_rs232_tx_stb <= 0;
    end
  end
  assign input_eth_rx_ack = s_input_eth_rx_ack;
  assign input_socket_ack = s_input_socket_ack;
  assign output_eth_tx_stb = s_output_eth_tx_stb;
  assign output_eth_tx = s_output_eth_tx;
  assign output_socket_stb = s_output_socket_stb;
  assign output_socket = s_output_socket;
  assign output_rs232_tx_stb = s_output_rs232_tx_stb;
  assign output_rs232_tx = s_output_rs232_tx;

endmodule
