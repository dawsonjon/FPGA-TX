//name : main_0
//input : input_eth_in:16
//output : output_audio_out:16
//output : output_eth_out:16
//source_file : /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c

///+============================================================================+
///|                                                                            |
///|                     This file was generated by Chips                       |
///|                                                                            |
///|                                  Chips                                     |
///|                                                                            |
///|                      http://github.com/dawsonjon/Chips-2.0                 |
///|                                                                            |
///|                                                             Python powered |
///+============================================================================+
module main_0(input_eth_in,input_eth_in_stb,output_audio_out_ack,output_eth_out_ack,clk,rst,output_audio_out,output_eth_out,output_audio_out_stb,output_eth_out_stb,input_eth_in_ack,exception);
  integer file_count;
  parameter  stop = 3'd0,
  instruction_fetch = 3'd1,
  operand_fetch = 3'd2,
  execute = 3'd3,
  load = 3'd4,
  wait_state = 3'd5,
  read = 3'd6,
  write = 3'd7;
  input [31:0] input_eth_in;
  input input_eth_in_stb;
  input output_audio_out_ack;
  input output_eth_out_ack;
  input clk;
  input rst;
  output [31:0] output_audio_out;
  output [31:0] output_eth_out;
  output output_audio_out_stb;
  output output_eth_out_stb;
  output input_eth_in_ack;
  reg [31:0] timer;
  reg [63:0] timer_clock;
  reg [15:0] program_counter;
  reg [15:0] program_counter_1;
  reg [15:0] program_counter_2;
  reg [44:0] instruction;
  reg [4:0] opcode_2;
  reg [3:0] a;
  reg [3:0] b;
  reg [3:0] z;
  reg write_enable;
  reg [3:0] address_a_2;
  reg [3:0] address_b_2;
  reg [3:0] address_z_2;
  reg [3:0] address_z_3;
  reg [31:0] load_data;
  reg [31:0] write_output;
  reg [31:0] write_value;
  reg [31:0] read_input;
  reg [15:0] literal_2;
  reg [31:0] a_hi;
  reg [31:0] b_hi;
  reg [31:0] a_lo;
  reg [31:0] b_lo;
  reg [63:0] long_result;
  reg [31:0] result;
  reg [15:0] address;
  reg [31:0] data_out;
  reg [31:0] data_in;
  reg [31:0] carry;
  reg [31:0] s_output_audio_out_stb;
  reg [31:0] s_output_eth_out_stb;
  reg [31:0] s_output_audio_out;
  reg [31:0] s_output_eth_out;
  reg [31:0] s_input_eth_in_ack;
  reg [7:0] state;
  output reg exception;
  reg [28:0] instructions [529:0];
  reg [31:0] memory [4096:0];
  reg [31:0] registers [15:0];
  wire [31:0] operand_a;
  wire [31:0] operand_b;
  wire [31:0] register_a;
  wire [31:0] register_b;
  wire [15:0] literal;
  wire [4:0] opcode;
  wire [3:0] address_a;
  wire [3:0] address_b;
  wire [3:0] address_z;
  wire [15:0] load_address;
  wire [15:0] store_address;
  wire [31:0] store_data;
  wire  store_enable;

  //////////////////////////////////////////////////////////////////////////////
  // INSTRUCTION INITIALIZATION                                                 
  //                                                                            
  // Initialise the contents of the instruction memory                          
  //
  // Intruction Set
  // ==============
  // 0 {'literal': True, 'op': 'literal'}
  // 1 {'literal': True, 'op': 'addl'}
  // 2 {'literal': False, 'op': 'store'}
  // 3 {'literal': True, 'op': 'call'}
  // 4 {'literal': False, 'op': 'stop'}
  // 5 {'literal': True, 'op': 'literal_hi'}
  // 6 {'literal': False, 'op': 'wait_clocks'}
  // 7 {'literal': False, 'op': 'load'}
  // 8 {'literal': False, 'op': 'unsigned_shift_right'}
  // 9 {'literal': False, 'op': 'unsigned_greater'}
  // 10 {'literal': True, 'op': 'jmp_if_false'}
  // 11 {'literal': False, 'op': 'add'}
  // 12 {'literal': False, 'op': 'write'}
  // 13 {'literal': True, 'op': 'goto'}
  // 14 {'literal': False, 'op': 'return'}
  // 15 {'literal': False, 'op': 'read'}
  // 16 {'literal': False, 'op': 'subtract'}
  // 17 {'literal': False, 'op': 'equal'}
  // Intructions
  // ===========
  
  initial
  begin
    instructions[0] = {5'd0, 4'd3, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 21 {'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 21, 'op': 'literal'}
    instructions[1] = {5'd0, 4'd4, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 21 {'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 21, 'op': 'literal'}
    instructions[2] = {5'd1, 4'd3, 4'd3, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 21 {'a': 3, 'literal': 10, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 21, 'op': 'addl'}
    instructions[3] = {5'd0, 4'd8, 4'd0, 16'd515};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 2 {'literal': 515, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 2, 'op': 'literal'}
    instructions[4] = {5'd0, 4'd2, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 2 {'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 2, 'op': 'literal'}
    instructions[5] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 2 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 2, 'op': 'store'}
    instructions[6] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 1 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 1, 'op': 'literal'}
    instructions[7] = {5'd0, 4'd2, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 1 {'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 1, 'op': 'literal'}
    instructions[8] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 1 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 1, 'op': 'store'}
    instructions[9] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 2 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 2, 'op': 'literal'}
    instructions[10] = {5'd0, 4'd2, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 2 {'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 2, 'op': 'literal'}
    instructions[11] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 2 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 2, 'op': 'store'}
    instructions[12] = {5'd0, 4'd8, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 4 {'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 4, 'op': 'literal'}
    instructions[13] = {5'd0, 4'd2, 4'd0, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 4 {'literal': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 4, 'op': 'literal'}
    instructions[14] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 4 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 4, 'op': 'store'}
    instructions[15] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 3 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 3, 'op': 'literal'}
    instructions[16] = {5'd0, 4'd2, 4'd0, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 3 {'literal': 7, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 3, 'op': 'literal'}
    instructions[17] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 3 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 3, 'op': 'store'}
    instructions[18] = {5'd0, 4'd8, 4'd0, 16'd1029};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 3 {'literal': 1029, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 3, 'op': 'literal'}
    instructions[19] = {5'd0, 4'd2, 4'd0, 16'd9};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 3 {'literal': 9, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 3, 'op': 'literal'}
    instructions[20] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 3 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 3, 'op': 'store'}
    instructions[21] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 21 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 21, 'op': 'addl'}
    instructions[22] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 21 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 21, 'op': 'addl'}
    instructions[23] = {5'd3, 4'd6, 4'd0, 16'd25};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 21 {'z': 6, 'label': 25, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 21, 'op': 'call'}
    instructions[24] = {5'd4, 4'd0, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 21 {'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 21, 'op': 'stop'}
    instructions[25] = {5'd1, 4'd3, 4'd3, 16'd258};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 7 {'a': 3, 'literal': 258, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 7, 'op': 'addl'}
    instructions[26] = {5'd0, 4'd8, 4'd0, 16'd61568};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 11 {'literal': 61568, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 11, 'op': 'literal'}
    instructions[27] = {5'd5, 4'd8, 4'd8, 16'd762};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 11 {'a': 8, 'literal': 762, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 11, 'op': 'literal_hi'}
    instructions[28] = {5'd6, 4'd0, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 11 {'a': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 11, 'op': 'wait_clocks'}
    instructions[29] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 14 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 14, 'op': 'store'}
    instructions[30] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 14 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 14, 'op': 'addl'}
    instructions[31] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 14 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 14, 'op': 'store'}
    instructions[32] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 14 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 14, 'op': 'addl'}
    instructions[33] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 14 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 14, 'op': 'addl'}
    instructions[34] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 14 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 14, 'op': 'store'}
    instructions[35] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 14 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 14, 'op': 'addl'}
    instructions[36] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 14 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 14, 'op': 'addl'}
    instructions[37] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 14 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 14, 'op': 'addl'}
    instructions[38] = {5'd3, 4'd6, 4'd0, 16'd133};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 14 {'z': 6, 'label': 133, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 14, 'op': 'call'}
    instructions[39] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 14 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 14, 'op': 'addl'}
    instructions[40] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 14 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 14, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[41] = {5'd7, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 14 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 14, 'op': 'load'}
    instructions[42] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 14 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 14, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[43] = {5'd7, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 14 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 14, 'op': 'load'}
    instructions[44] = {5'd0, 4'd2, 4'd0, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 14 {'literal': 4, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 14, 'op': 'literal'}
    instructions[45] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 14 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 14, 'op': 'load'}
    instructions[46] = {5'd1, 4'd2, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 14 {'a': 4, 'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 14, 'op': 'addl'}
    instructions[47] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 14 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 14, 'op': 'store'}
    instructions[48] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 15 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 15, 'op': 'store'}
    instructions[49] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 15 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 15, 'op': 'addl'}
    instructions[50] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 15 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 15, 'op': 'store'}
    instructions[51] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 15 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 15, 'op': 'addl'}
    instructions[52] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 15 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 15, 'op': 'addl'}
    instructions[53] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 15 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 15, 'op': 'store'}
    instructions[54] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 15 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 15, 'op': 'addl'}
    instructions[55] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 15 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 15, 'op': 'addl'}
    instructions[56] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 15 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 15, 'op': 'addl'}
    instructions[57] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 15 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 15, 'op': 'load'}
    instructions[58] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 15 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 15, 'op': 'store'}
    instructions[59] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 15 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 15, 'op': 'addl'}
    instructions[60] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 15 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 15, 'op': 'addl'}
    instructions[61] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 15 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 15, 'op': 'addl'}
    instructions[62] = {5'd3, 4'd6, 4'd0, 16'd343};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 15 {'z': 6, 'label': 343, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 15, 'op': 'call'}
    instructions[63] = {5'd1, 4'd3, 4'd3, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 15 {'a': 3, 'literal': -2, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 15, 'op': 'addl'}
    instructions[64] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 15 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 15, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[65] = {5'd7, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 15 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 15, 'op': 'load'}
    instructions[66] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 15 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 15, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[67] = {5'd7, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 15 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 15, 'op': 'load'}
    instructions[68] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 15 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 15, 'op': 'addl'}
    instructions[69] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16, 'op': 'literal'}
    instructions[70] = {5'd1, 4'd2, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16, 'op': 'addl'}
    instructions[71] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16, 'op': 'store'}
    instructions[72] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16, 'op': 'addl'}
    instructions[73] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16, 'op': 'addl'}
    instructions[74] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16, 'op': 'load'}
    instructions[75] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16, 'op': 'store'}
    instructions[76] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16, 'op': 'addl'}
    instructions[77] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16, 'op': 'literal'}
    instructions[78] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16, 'op': 'store'}
    instructions[79] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16, 'op': 'addl'}
    instructions[80] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16, 'op': 'addl'}
    instructions[81] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16, 'op': 'addl'}
    instructions[82] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16, 'op': 'load'}
    instructions[83] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[84] = {5'd7, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16, 'op': 'load'}
    instructions[85] = {5'd8, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16, 'op': 'unsigned_shift_right'}
    instructions[86] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[87] = {5'd7, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16, 'op': 'load'}
    instructions[88] = {5'd9, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16, 'op': 'unsigned_greater'}
    instructions[89] = {5'd10, 4'd0, 4'd8, 16'd129};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16 {'a': 8, 'label': 129, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16, 'op': 'jmp_if_false'}
    instructions[90] = {5'd0, 4'd8, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 17 {'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 17, 'op': 'literal'}
    instructions[91] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 17 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 17, 'op': 'addl'}
    instructions[92] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 17 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 17, 'op': 'load'}
    instructions[93] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 17 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 17, 'op': 'store'}
    instructions[94] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 17 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 17, 'op': 'addl'}
    instructions[95] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 17 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 17, 'op': 'addl'}
    instructions[96] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 17 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 17, 'op': 'store'}
    instructions[97] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 17 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 17, 'op': 'addl'}
    instructions[98] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 17 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 17, 'op': 'addl'}
    instructions[99] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 17 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 17, 'op': 'addl'}
    instructions[100] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 17 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 17, 'op': 'load'}
    instructions[101] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 17 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 17, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[102] = {5'd7, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 17 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 17, 'op': 'load'}
    instructions[103] = {5'd11, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 17 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 17, 'op': 'add'}
    instructions[104] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 17 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 17, 'op': 'addl'}
    instructions[105] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 17 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 17, 'op': 'load'}
    instructions[106] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 17 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 17, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[107] = {5'd7, 4'd0, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 17 {'a': 3, 'z': 0, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 17, 'op': 'load'}
    instructions[108] = {5'd12, 4'd0, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 17 {'a': 0, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 17, 'op': 'write'}
    instructions[109] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 17 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 17, 'op': 'addl'}
    instructions[110] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16, 'op': 'addl'}
    instructions[111] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16, 'op': 'addl'}
    instructions[112] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16, 'op': 'load'}
    instructions[113] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16, 'op': 'store'}
    instructions[114] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16, 'op': 'addl'}
    instructions[115] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16, 'op': 'literal'}
    instructions[116] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16, 'op': 'store'}
    instructions[117] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16, 'op': 'addl'}
    instructions[118] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16, 'op': 'addl'}
    instructions[119] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16, 'op': 'addl'}
    instructions[120] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16, 'op': 'load'}
    instructions[121] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[122] = {5'd7, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16, 'op': 'load'}
    instructions[123] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16, 'op': 'add'}
    instructions[124] = {5'd1, 4'd2, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16, 'op': 'addl'}
    instructions[125] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16, 'op': 'store'}
    instructions[126] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[127] = {5'd7, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16, 'op': 'load'}
    instructions[128] = {5'd13, 4'd0, 4'd0, 16'd72};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16 {'label': 72, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 16, 'op': 'goto'}
    instructions[129] = {5'd13, 4'd0, 4'd0, 16'd29};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 13 {'label': 29, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 13, 'op': 'goto'}
    instructions[130] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 7 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 7, 'op': 'addl'}
    instructions[131] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 7 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 7, 'op': 'addl'}
    instructions[132] = {5'd14, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 7 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/application.c : 7, 'op': 'return'}
    instructions[133] = {5'd1, 4'd3, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 7 {'a': 3, 'literal': 8, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 7, 'op': 'addl'}
    instructions[134] = {5'd0, 4'd8, 4'd0, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 13 {'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 13, 'op': 'literal'}
    instructions[135] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 13 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 13, 'op': 'addl'}
    instructions[136] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 13 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 13, 'op': 'load'}
    instructions[137] = {5'd15, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 13 {'a': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 13, 'op': 'read'}
    instructions[138] = {5'd1, 4'd2, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 13 {'a': 4, 'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 13, 'op': 'addl'}
    instructions[139] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 13 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 13, 'op': 'store'}
    instructions[140] = {5'd0, 4'd8, 4'd0, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 14 {'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 14, 'op': 'literal'}
    instructions[141] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 14 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 14, 'op': 'addl'}
    instructions[142] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 14 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 14, 'op': 'load'}
    instructions[143] = {5'd15, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 14 {'a': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 14, 'op': 'read'}
    instructions[144] = {5'd1, 4'd2, 4'd4, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 14 {'a': 4, 'literal': 4, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 14, 'op': 'addl'}
    instructions[145] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 14 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 14, 'op': 'store'}
    instructions[146] = {5'd0, 4'd8, 4'd0, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 15 {'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 15, 'op': 'literal'}
    instructions[147] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 15 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 15, 'op': 'addl'}
    instructions[148] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 15 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 15, 'op': 'load'}
    instructions[149] = {5'd15, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 15 {'a': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 15, 'op': 'read'}
    instructions[150] = {5'd1, 4'd2, 4'd4, 16'd5};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 15 {'a': 4, 'literal': 5, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 15, 'op': 'addl'}
    instructions[151] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 15 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 15, 'op': 'store'}
    instructions[152] = {5'd0, 4'd8, 4'd0, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 16 {'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 16, 'op': 'literal'}
    instructions[153] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 16 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 16, 'op': 'addl'}
    instructions[154] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 16 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 16, 'op': 'load'}
    instructions[155] = {5'd15, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 16 {'a': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 16, 'op': 'read'}
    instructions[156] = {5'd1, 4'd2, 4'd4, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 16 {'a': 4, 'literal': 6, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 16, 'op': 'addl'}
    instructions[157] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 16 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 16, 'op': 'store'}
    instructions[158] = {5'd0, 4'd8, 4'd0, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 17 {'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 17, 'op': 'literal'}
    instructions[159] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 17 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 17, 'op': 'addl'}
    instructions[160] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 17 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 17, 'op': 'load'}
    instructions[161] = {5'd15, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 17 {'a': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 17, 'op': 'read'}
    instructions[162] = {5'd0, 4'd2, 4'd0, 16'd5};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 17 {'literal': 5, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 17, 'op': 'literal'}
    instructions[163] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 17 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 17, 'op': 'store'}
    instructions[164] = {5'd0, 4'd8, 4'd0, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 18 {'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 18, 'op': 'literal'}
    instructions[165] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 18 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 18, 'op': 'addl'}
    instructions[166] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 18 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 18, 'op': 'load'}
    instructions[167] = {5'd15, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 18 {'a': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 18, 'op': 'read'}
    instructions[168] = {5'd0, 4'd2, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 18 {'literal': 8, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 18, 'op': 'literal'}
    instructions[169] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 18 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 18, 'op': 'store'}
    instructions[170] = {5'd0, 4'd8, 4'd0, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 19 {'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 19, 'op': 'literal'}
    instructions[171] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 19 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 19, 'op': 'addl'}
    instructions[172] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 19 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 19, 'op': 'load'}
    instructions[173] = {5'd15, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 19 {'a': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 19, 'op': 'read'}
    instructions[174] = {5'd0, 4'd2, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 19 {'literal': 6, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 19, 'op': 'literal'}
    instructions[175] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 19 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 19, 'op': 'store'}
    instructions[176] = {5'd0, 4'd8, 4'd0, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 20 {'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 20, 'op': 'literal'}
    instructions[177] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 20 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 20, 'op': 'addl'}
    instructions[178] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 20 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 20, 'op': 'load'}
    instructions[179] = {5'd15, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 20 {'a': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 20, 'op': 'read'}
    instructions[180] = {5'd1, 4'd2, 4'd4, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 20 {'a': 4, 'literal': 7, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 20, 'op': 'addl'}
    instructions[181] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 20 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 20, 'op': 'store'}
    instructions[182] = {5'd0, 4'd8, 4'd0, 16'd14};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 21 {'literal': 14, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 21, 'op': 'literal'}
    instructions[183] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 21 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 21, 'op': 'store'}
    instructions[184] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 21 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 21, 'op': 'addl'}
    instructions[185] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 21 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 21, 'op': 'addl'}
    instructions[186] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 21 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 21, 'op': 'addl'}
    instructions[187] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 21 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 21, 'op': 'load'}
    instructions[188] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 21 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 21, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[189] = {5'd7, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 21 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 21, 'op': 'load'}
    instructions[190] = {5'd16, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 21 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 21, 'op': 'subtract'}
    instructions[191] = {5'd1, 4'd2, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 21 {'a': 4, 'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 21, 'op': 'addl'}
    instructions[192] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 21 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 21, 'op': 'store'}
    instructions[193] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 22 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 22, 'op': 'literal'}
    instructions[194] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 22 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 22, 'op': 'store'}
    instructions[195] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 22 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 22, 'op': 'addl'}
    instructions[196] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 22 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 22, 'op': 'literal'}
    instructions[197] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 22 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 22, 'op': 'store'}
    instructions[198] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 22 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 22, 'op': 'addl'}
    instructions[199] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 22 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 22, 'op': 'addl'}
    instructions[200] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 22 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 22, 'op': 'addl'}
    instructions[201] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 22 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 22, 'op': 'load'}
    instructions[202] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 22 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 22, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[203] = {5'd7, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 22 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 22, 'op': 'load'}
    instructions[204] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 22 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 22, 'op': 'add'}
    instructions[205] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 22 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 22, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[206] = {5'd7, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 22 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 22, 'op': 'load'}
    instructions[207] = {5'd8, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 22 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 22, 'op': 'unsigned_shift_right'}
    instructions[208] = {5'd1, 4'd2, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 22 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 22, 'op': 'addl'}
    instructions[209] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 22 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 22, 'op': 'store'}
    instructions[210] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24, 'op': 'literal'}
    instructions[211] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24, 'op': 'store'}
    instructions[212] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24, 'op': 'addl'}
    instructions[213] = {5'd1, 4'd8, 4'd4, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24 {'a': 4, 'literal': 4, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24, 'op': 'addl'}
    instructions[214] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24, 'op': 'addl'}
    instructions[215] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24, 'op': 'load'}
    instructions[216] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[217] = {5'd7, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24, 'op': 'load'}
    instructions[218] = {5'd17, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24, 'op': 'equal'}
    instructions[219] = {5'd10, 4'd0, 4'd8, 16'd229};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24 {'a': 8, 'label': 229, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24, 'op': 'jmp_if_false'}
    instructions[220] = {5'd0, 4'd8, 4'd0, 16'd515};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24 {'literal': 515, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24, 'op': 'literal'}
    instructions[221] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24, 'op': 'store'}
    instructions[222] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24, 'op': 'addl'}
    instructions[223] = {5'd1, 4'd8, 4'd4, 16'd5};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24 {'a': 4, 'literal': 5, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24, 'op': 'addl'}
    instructions[224] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24, 'op': 'addl'}
    instructions[225] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24, 'op': 'load'}
    instructions[226] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[227] = {5'd7, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24, 'op': 'load'}
    instructions[228] = {5'd17, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24, 'op': 'equal'}
    instructions[229] = {5'd10, 4'd0, 4'd8, 16'd239};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24 {'a': 8, 'label': 239, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24, 'op': 'jmp_if_false'}
    instructions[230] = {5'd0, 4'd8, 4'd0, 16'd1029};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24 {'literal': 1029, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24, 'op': 'literal'}
    instructions[231] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24, 'op': 'store'}
    instructions[232] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24, 'op': 'addl'}
    instructions[233] = {5'd1, 4'd8, 4'd4, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24 {'a': 4, 'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24, 'op': 'addl'}
    instructions[234] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24, 'op': 'addl'}
    instructions[235] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24, 'op': 'load'}
    instructions[236] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[237] = {5'd7, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24, 'op': 'load'}
    instructions[238] = {5'd17, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24, 'op': 'equal'}
    instructions[239] = {5'd10, 4'd0, 4'd8, 16'd313};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24 {'a': 8, 'label': 313, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24, 'op': 'jmp_if_false'}
    instructions[240] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 26 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 26, 'op': 'literal'}
    instructions[241] = {5'd1, 4'd2, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 26 {'a': 4, 'literal': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 26, 'op': 'addl'}
    instructions[242] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 26 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 26, 'op': 'store'}
    instructions[243] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 27 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 27, 'op': 'addl'}
    instructions[244] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 27 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 27, 'op': 'addl'}
    instructions[245] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 27 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 27, 'op': 'load'}
    instructions[246] = {5'd10, 4'd0, 4'd8, 16'd302};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 31 {'a': 8, 'label': 302, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 31, 'op': 'jmp_if_false'}
    instructions[247] = {5'd0, 4'd8, 4'd0, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28 {'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28, 'op': 'literal'}
    instructions[248] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28, 'op': 'addl'}
    instructions[249] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28, 'op': 'load'}
    instructions[250] = {5'd15, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28 {'a': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28, 'op': 'read'}
    instructions[251] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28, 'op': 'store'}
    instructions[252] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28, 'op': 'addl'}
    instructions[253] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28, 'op': 'addl'}
    instructions[254] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28, 'op': 'addl'}
    instructions[255] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28, 'op': 'load'}
    instructions[256] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28, 'op': 'store'}
    instructions[257] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28, 'op': 'addl'}
    instructions[258] = {5'd1, 4'd8, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28 {'a': 4, 'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28, 'op': 'addl'}
    instructions[259] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28, 'op': 'addl'}
    instructions[260] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28, 'op': 'load'}
    instructions[261] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28, 'op': 'store'}
    instructions[262] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28, 'op': 'addl'}
    instructions[263] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28, 'op': 'literal'}
    instructions[264] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28, 'op': 'store'}
    instructions[265] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28, 'op': 'addl'}
    instructions[266] = {5'd1, 4'd8, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28 {'a': 4, 'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28, 'op': 'addl'}
    instructions[267] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28, 'op': 'addl'}
    instructions[268] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28, 'op': 'load'}
    instructions[269] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[270] = {5'd7, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28, 'op': 'load'}
    instructions[271] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28, 'op': 'add'}
    instructions[272] = {5'd1, 4'd2, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28 {'a': 4, 'literal': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28, 'op': 'addl'}
    instructions[273] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28, 'op': 'store'}
    instructions[274] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[275] = {5'd7, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28, 'op': 'load'}
    instructions[276] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[277] = {5'd7, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28, 'op': 'load'}
    instructions[278] = {5'd11, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28, 'op': 'add'}
    instructions[279] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28, 'op': 'addl'}
    instructions[280] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[281] = {5'd7, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28, 'op': 'load'}
    instructions[282] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 28, 'op': 'store'}
    instructions[283] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 29 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 29, 'op': 'addl'}
    instructions[284] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 29 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 29, 'op': 'addl'}
    instructions[285] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 29 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 29, 'op': 'load'}
    instructions[286] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 29 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 29, 'op': 'store'}
    instructions[287] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 29 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 29, 'op': 'addl'}
    instructions[288] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 29 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 29, 'op': 'literal'}
    instructions[289] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 29 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 29, 'op': 'store'}
    instructions[290] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 29 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 29, 'op': 'addl'}
    instructions[291] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 29 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 29, 'op': 'addl'}
    instructions[292] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 29 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 29, 'op': 'addl'}
    instructions[293] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 29 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 29, 'op': 'load'}
    instructions[294] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 29 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 29, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[295] = {5'd7, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 29 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 29, 'op': 'load'}
    instructions[296] = {5'd16, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 29 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 29, 'op': 'subtract'}
    instructions[297] = {5'd1, 4'd2, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 29 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 29, 'op': 'addl'}
    instructions[298] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 29 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 29, 'op': 'store'}
    instructions[299] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 29 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 29, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[300] = {5'd7, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 29 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 29, 'op': 'load'}
    instructions[301] = {5'd13, 4'd0, 4'd0, 16'd303};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 31 {'label': 303, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 31, 'op': 'goto'}
    instructions[302] = {5'd13, 4'd0, 4'd0, 16'd304};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 31 {'label': 304, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 31, 'op': 'goto'}
    instructions[303] = {5'd13, 4'd0, 4'd0, 16'd243};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 27 {'label': 243, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 27, 'op': 'goto'}
    instructions[304] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 31 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 31, 'op': 'addl'}
    instructions[305] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 31 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 31, 'op': 'addl'}
    instructions[306] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 31 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 31, 'op': 'load'}
    instructions[307] = {5'd0, 4'd2, 4'd0, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 31 {'literal': 4, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 31, 'op': 'literal'}
    instructions[308] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 31 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 31, 'op': 'store'}
    instructions[309] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 31 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 31, 'op': 'addl'}
    instructions[310] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 31 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 31, 'op': 'addl'}
    instructions[311] = {5'd14, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 31 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 31, 'op': 'return'}
    instructions[312] = {5'd13, 4'd0, 4'd0, 16'd342};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24 {'label': 342, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 24, 'op': 'goto'}
    instructions[313] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 35 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 35, 'op': 'addl'}
    instructions[314] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 35 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 35, 'op': 'addl'}
    instructions[315] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 35 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 35, 'op': 'load'}
    instructions[316] = {5'd10, 4'd0, 4'd8, 16'd340};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 40 {'a': 8, 'label': 340, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 40, 'op': 'jmp_if_false'}
    instructions[317] = {5'd0, 4'd8, 4'd0, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 36 {'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 36, 'op': 'literal'}
    instructions[318] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 36 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 36, 'op': 'addl'}
    instructions[319] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 36 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 36, 'op': 'load'}
    instructions[320] = {5'd15, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 36 {'a': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 36, 'op': 'read'}
    instructions[321] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 37 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 37, 'op': 'addl'}
    instructions[322] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 37 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 37, 'op': 'addl'}
    instructions[323] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 37 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 37, 'op': 'load'}
    instructions[324] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 37 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 37, 'op': 'store'}
    instructions[325] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 37 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 37, 'op': 'addl'}
    instructions[326] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 37 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 37, 'op': 'literal'}
    instructions[327] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 37 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 37, 'op': 'store'}
    instructions[328] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 37 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 37, 'op': 'addl'}
    instructions[329] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 37 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 37, 'op': 'addl'}
    instructions[330] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 37 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 37, 'op': 'addl'}
    instructions[331] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 37 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 37, 'op': 'load'}
    instructions[332] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 37 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 37, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[333] = {5'd7, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 37 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 37, 'op': 'load'}
    instructions[334] = {5'd16, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 37 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 37, 'op': 'subtract'}
    instructions[335] = {5'd1, 4'd2, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 37 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 37, 'op': 'addl'}
    instructions[336] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 37 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 37, 'op': 'store'}
    instructions[337] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 37 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 37, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[338] = {5'd7, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 37 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 37, 'op': 'load'}
    instructions[339] = {5'd13, 4'd0, 4'd0, 16'd341};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 40 {'label': 341, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 40, 'op': 'goto'}
    instructions[340] = {5'd13, 4'd0, 4'd0, 16'd342};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 40 {'label': 342, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 40, 'op': 'goto'}
    instructions[341] = {5'd13, 4'd0, 4'd0, 16'd313};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 35 {'label': 313, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 35, 'op': 'goto'}
    instructions[342] = {5'd13, 4'd0, 4'd0, 16'd134};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 12 {'label': 134, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 12, 'op': 'goto'}
    instructions[343] = {5'd1, 4'd3, 4'd3, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 45 {'a': 3, 'literal': 3, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 45, 'op': 'addl'}
    instructions[344] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 49 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 49, 'op': 'literal'}
    instructions[345] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 49 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 49, 'op': 'store'}
    instructions[346] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 49 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 49, 'op': 'addl'}
    instructions[347] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 49 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 49, 'op': 'literal'}
    instructions[348] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 49 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 49, 'op': 'store'}
    instructions[349] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 49 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 49, 'op': 'addl'}
    instructions[350] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 49 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 49, 'op': 'addl'}
    instructions[351] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 49 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 49, 'op': 'addl'}
    instructions[352] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 49 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 49, 'op': 'load'}
    instructions[353] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 49 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 49, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[354] = {5'd7, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 49 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 49, 'op': 'load'}
    instructions[355] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 49 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 49, 'op': 'add'}
    instructions[356] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 49 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 49, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[357] = {5'd7, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 49 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 49, 'op': 'load'}
    instructions[358] = {5'd8, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 49 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 49, 'op': 'unsigned_shift_right'}
    instructions[359] = {5'd1, 4'd2, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 49 {'a': 4, 'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 49, 'op': 'addl'}
    instructions[360] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 49 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 49, 'op': 'store'}
    instructions[361] = {5'd0, 4'd8, 4'd0, 16'd14};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 50 {'literal': 14, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 50, 'op': 'literal'}
    instructions[362] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 50 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 50, 'op': 'store'}
    instructions[363] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 50 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 50, 'op': 'addl'}
    instructions[364] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 50 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 50, 'op': 'addl'}
    instructions[365] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 50 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 50, 'op': 'addl'}
    instructions[366] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 50 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 50, 'op': 'load'}
    instructions[367] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 50 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 50, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[368] = {5'd7, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 50 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 50, 'op': 'load'}
    instructions[369] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 50 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 50, 'op': 'add'}
    instructions[370] = {5'd1, 4'd2, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 50 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 50, 'op': 'addl'}
    instructions[371] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 50 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 50, 'op': 'store'}
    instructions[372] = {5'd0, 4'd8, 4'd0, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 52 {'literal': 7, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 52, 'op': 'literal'}
    instructions[373] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 52 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 52, 'op': 'addl'}
    instructions[374] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 52 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 52, 'op': 'load'}
    instructions[375] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 52 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 52, 'op': 'store'}
    instructions[376] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 52 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 52, 'op': 'addl'}
    instructions[377] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 52 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 52, 'op': 'addl'}
    instructions[378] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 52 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 52, 'op': 'addl'}
    instructions[379] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 52 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 52, 'op': 'load'}
    instructions[380] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 52 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 52, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[381] = {5'd7, 4'd0, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 52 {'a': 3, 'z': 0, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 52, 'op': 'load'}
    instructions[382] = {5'd12, 4'd0, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 52 {'a': 0, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 52, 'op': 'write'}
    instructions[383] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 52 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 52, 'op': 'addl'}
    instructions[384] = {5'd0, 4'd8, 4'd0, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 53 {'literal': 7, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 53, 'op': 'literal'}
    instructions[385] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 53 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 53, 'op': 'addl'}
    instructions[386] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 53 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 53, 'op': 'load'}
    instructions[387] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 53 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 53, 'op': 'store'}
    instructions[388] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 53 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 53, 'op': 'addl'}
    instructions[389] = {5'd0, 4'd8, 4'd0, 16'd5};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 53 {'literal': 5, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 53, 'op': 'literal'}
    instructions[390] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 53 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 53, 'op': 'addl'}
    instructions[391] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 53 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 53, 'op': 'load'}
    instructions[392] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 53 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 53, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[393] = {5'd7, 4'd0, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 53 {'a': 3, 'z': 0, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 53, 'op': 'load'}
    instructions[394] = {5'd12, 4'd0, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 53 {'a': 0, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 53, 'op': 'write'}
    instructions[395] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 53 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 53, 'op': 'addl'}
    instructions[396] = {5'd0, 4'd8, 4'd0, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 54 {'literal': 7, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 54, 'op': 'literal'}
    instructions[397] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 54 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 54, 'op': 'addl'}
    instructions[398] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 54 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 54, 'op': 'load'}
    instructions[399] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 54 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 54, 'op': 'store'}
    instructions[400] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 54 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 54, 'op': 'addl'}
    instructions[401] = {5'd0, 4'd8, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 54 {'literal': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 54, 'op': 'literal'}
    instructions[402] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 54 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 54, 'op': 'addl'}
    instructions[403] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 54 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 54, 'op': 'load'}
    instructions[404] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 54 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 54, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[405] = {5'd7, 4'd0, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 54 {'a': 3, 'z': 0, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 54, 'op': 'load'}
    instructions[406] = {5'd12, 4'd0, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 54 {'a': 0, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 54, 'op': 'write'}
    instructions[407] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 54 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 54, 'op': 'addl'}
    instructions[408] = {5'd0, 4'd8, 4'd0, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 55 {'literal': 7, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 55, 'op': 'literal'}
    instructions[409] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 55 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 55, 'op': 'addl'}
    instructions[410] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 55 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 55, 'op': 'load'}
    instructions[411] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 55 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 55, 'op': 'store'}
    instructions[412] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 55 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 55, 'op': 'addl'}
    instructions[413] = {5'd0, 4'd8, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 55 {'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 55, 'op': 'literal'}
    instructions[414] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 55 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 55, 'op': 'addl'}
    instructions[415] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 55 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 55, 'op': 'load'}
    instructions[416] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 55 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 55, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[417] = {5'd7, 4'd0, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 55 {'a': 3, 'z': 0, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 55, 'op': 'load'}
    instructions[418] = {5'd12, 4'd0, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 55 {'a': 0, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 55, 'op': 'write'}
    instructions[419] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 55 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 55, 'op': 'addl'}
    instructions[420] = {5'd0, 4'd8, 4'd0, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 56 {'literal': 7, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 56, 'op': 'literal'}
    instructions[421] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 56 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 56, 'op': 'addl'}
    instructions[422] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 56 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 56, 'op': 'load'}
    instructions[423] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 56 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 56, 'op': 'store'}
    instructions[424] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 56 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 56, 'op': 'addl'}
    instructions[425] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 56 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 56, 'op': 'literal'}
    instructions[426] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 56 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 56, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[427] = {5'd7, 4'd0, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 56 {'a': 3, 'z': 0, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 56, 'op': 'load'}
    instructions[428] = {5'd12, 4'd0, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 56 {'a': 0, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 56, 'op': 'write'}
    instructions[429] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 56 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 56, 'op': 'addl'}
    instructions[430] = {5'd0, 4'd8, 4'd0, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 57 {'literal': 7, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 57, 'op': 'literal'}
    instructions[431] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 57 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 57, 'op': 'addl'}
    instructions[432] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 57 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 57, 'op': 'load'}
    instructions[433] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 57 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 57, 'op': 'store'}
    instructions[434] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 57 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 57, 'op': 'addl'}
    instructions[435] = {5'd0, 4'd8, 4'd0, 16'd515};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 57 {'literal': 515, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 57, 'op': 'literal'}
    instructions[436] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 57 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 57, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[437] = {5'd7, 4'd0, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 57 {'a': 3, 'z': 0, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 57, 'op': 'load'}
    instructions[438] = {5'd12, 4'd0, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 57 {'a': 0, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 57, 'op': 'write'}
    instructions[439] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 57 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 57, 'op': 'addl'}
    instructions[440] = {5'd0, 4'd8, 4'd0, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 58 {'literal': 7, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 58, 'op': 'literal'}
    instructions[441] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 58 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 58, 'op': 'addl'}
    instructions[442] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 58 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 58, 'op': 'load'}
    instructions[443] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 58 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 58, 'op': 'store'}
    instructions[444] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 58 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 58, 'op': 'addl'}
    instructions[445] = {5'd0, 4'd8, 4'd0, 16'd1029};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 58 {'literal': 1029, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 58, 'op': 'literal'}
    instructions[446] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 58 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 58, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[447] = {5'd7, 4'd0, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 58 {'a': 3, 'z': 0, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 58, 'op': 'load'}
    instructions[448] = {5'd12, 4'd0, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 58 {'a': 0, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 58, 'op': 'write'}
    instructions[449] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 58 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 58, 'op': 'addl'}
    instructions[450] = {5'd0, 4'd8, 4'd0, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 59 {'literal': 7, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 59, 'op': 'literal'}
    instructions[451] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 59 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 59, 'op': 'addl'}
    instructions[452] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 59 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 59, 'op': 'load'}
    instructions[453] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 59 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 59, 'op': 'store'}
    instructions[454] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 59 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 59, 'op': 'addl'}
    instructions[455] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 59 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 59, 'op': 'addl'}
    instructions[456] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 59 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 59, 'op': 'addl'}
    instructions[457] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 59 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 59, 'op': 'load'}
    instructions[458] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 59 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 59, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[459] = {5'd7, 4'd0, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 59 {'a': 3, 'z': 0, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 59, 'op': 'load'}
    instructions[460] = {5'd12, 4'd0, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 59 {'a': 0, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 59, 'op': 'write'}
    instructions[461] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 59 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 59, 'op': 'addl'}
    instructions[462] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 61 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 61, 'op': 'literal'}
    instructions[463] = {5'd1, 4'd2, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 61 {'a': 4, 'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 61, 'op': 'addl'}
    instructions[464] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 61 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 61, 'op': 'store'}
    instructions[465] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 62 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 62, 'op': 'addl'}
    instructions[466] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 62 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 62, 'op': 'addl'}
    instructions[467] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 62 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 62, 'op': 'load'}
    instructions[468] = {5'd10, 4'd0, 4'd8, 16'd525};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 67 {'a': 8, 'label': 525, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 67, 'op': 'jmp_if_false'}
    instructions[469] = {5'd0, 4'd8, 4'd0, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63 {'literal': 7, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63, 'op': 'literal'}
    instructions[470] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63, 'op': 'addl'}
    instructions[471] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63, 'op': 'load'}
    instructions[472] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63, 'op': 'store'}
    instructions[473] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63, 'op': 'addl'}
    instructions[474] = {5'd1, 4'd8, 4'd4, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63 {'a': 4, 'literal': -2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63, 'op': 'addl'}
    instructions[475] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63, 'op': 'addl'}
    instructions[476] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63, 'op': 'load'}
    instructions[477] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63, 'op': 'store'}
    instructions[478] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63, 'op': 'addl'}
    instructions[479] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63, 'op': 'addl'}
    instructions[480] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63, 'op': 'addl'}
    instructions[481] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63, 'op': 'load'}
    instructions[482] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63, 'op': 'store'}
    instructions[483] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63, 'op': 'addl'}
    instructions[484] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63, 'op': 'literal'}
    instructions[485] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63, 'op': 'store'}
    instructions[486] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63, 'op': 'addl'}
    instructions[487] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63, 'op': 'addl'}
    instructions[488] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63, 'op': 'addl'}
    instructions[489] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63, 'op': 'load'}
    instructions[490] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[491] = {5'd7, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63, 'op': 'load'}
    instructions[492] = {5'd11, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63, 'op': 'add'}
    instructions[493] = {5'd1, 4'd2, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63 {'a': 4, 'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63, 'op': 'addl'}
    instructions[494] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63, 'op': 'store'}
    instructions[495] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[496] = {5'd7, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63, 'op': 'load'}
    instructions[497] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[498] = {5'd7, 4'd2, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63 {'a': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63, 'op': 'load'}
    instructions[499] = {5'd11, 4'd8, 4'd8, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63 {'a': 8, 'z': 8, 'b': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63, 'op': 'add'}
    instructions[500] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63, 'op': 'addl'}
    instructions[501] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63, 'op': 'load'}
    instructions[502] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[503] = {5'd7, 4'd0, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63 {'a': 3, 'z': 0, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63, 'op': 'load'}
    instructions[504] = {5'd12, 4'd0, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63 {'a': 0, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63, 'op': 'write'}
    instructions[505] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 63, 'op': 'addl'}
    instructions[506] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 64 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 64, 'op': 'addl'}
    instructions[507] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 64 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 64, 'op': 'addl'}
    instructions[508] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 64 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 64, 'op': 'load'}
    instructions[509] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 64 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 64, 'op': 'store'}
    instructions[510] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 64 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 64, 'op': 'addl'}
    instructions[511] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 64 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 64, 'op': 'literal'}
    instructions[512] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 64 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 64, 'op': 'store'}
    instructions[513] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 64 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 64, 'op': 'addl'}
    instructions[514] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 64 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 64, 'op': 'addl'}
    instructions[515] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 64 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 64, 'op': 'addl'}
    instructions[516] = {5'd7, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 64 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 64, 'op': 'load'}
    instructions[517] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 64 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 64, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[518] = {5'd7, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 64 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 64, 'op': 'load'}
    instructions[519] = {5'd16, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 64 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 64, 'op': 'subtract'}
    instructions[520] = {5'd1, 4'd2, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 64 {'a': 4, 'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 64, 'op': 'addl'}
    instructions[521] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 64 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 64, 'op': 'store'}
    instructions[522] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 64 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 64, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[523] = {5'd7, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 64 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 64, 'op': 'load'}
    instructions[524] = {5'd13, 4'd0, 4'd0, 16'd526};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 67 {'label': 526, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 67, 'op': 'goto'}
    instructions[525] = {5'd13, 4'd0, 4'd0, 16'd527};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 67 {'label': 527, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 67, 'op': 'goto'}
    instructions[526] = {5'd13, 4'd0, 4'd0, 16'd465};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 62 {'label': 465, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 62, 'op': 'goto'}
    instructions[527] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 45 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 45, 'op': 'addl'}
    instructions[528] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 45 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 45, 'op': 'addl'}
    instructions[529] = {5'd14, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 45 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/audio_output/ethernet.h : 45, 'op': 'return'}
  end

  
  always @(posedge clk)
  begin
    load_data <= memory[load_address];
    if(store_enable && state == execute) begin
      memory[store_address] <= store_data;
    end
  end


  //////////////////////////////////////////////////////////////////////////////
  // PIPELINE STAGE 1 -- FETCH INSTRUCTION
  //                                                                            
  
  always @(posedge clk)
  begin
    //implement memory for instructions
    if (state == instruction_fetch || state == operand_fetch || state == execute) begin
      instruction <= instructions[program_counter];
      program_counter_1 <= program_counter;
    end
  end

  assign opcode    = instruction[28:24];
  assign address_z = instruction[23:20];
  assign address_a = instruction[19:16];
  assign address_b = instruction[3:0];
  assign literal   = instruction[15:0];

  //////////////////////////////////////////////////////////////////////////////
  // PIPELINE STAGE 2 -- FETCH OPERANDS
  //                                                                            
  
  always @(posedge clk)
  begin
    if (write_enable) begin
      registers[address_z_3] <= result;
    end
    if (state == operand_fetch || state == execute) begin
      opcode_2 <= opcode;
      literal_2 <= literal;
      address_a_2 <= address_a;
      address_b_2 <= address_b;
      address_z_2 <= address_z;
      program_counter_2 <= program_counter_1;
    end
  end
  assign register_a = registers[address_a_2];
  assign register_b = registers[address_b_2];
  assign operand_a = (address_a_2 == address_z_3 && write_enable)?result:register_a;
  assign operand_b = (address_b_2 == address_z_3 && write_enable)?result:register_b;
  assign store_address = operand_a;
  assign load_address = operand_a;
  assign store_data = operand_b;
  assign store_enable = (opcode_2==2);

  //////////////////////////////////////////////////////////////////////////////
  // PIPELINE STAGE 3 -- EXECUTE
  //                                                                            
  
  always @(posedge clk)
  begin

  write_enable <= 0;
  timer_clock <= timer_clock + 1;
  case(state)

    //instruction_fetch
    instruction_fetch: begin
      program_counter <= program_counter + 1;
      state <= operand_fetch;
    end
    //operand_fetch
    operand_fetch: begin
      program_counter <= program_counter + 1;
      state <= execute;
    end
    //execute
    execute: begin
      program_counter <= program_counter + 1;
      address_z_3 <= address_z_2;
      case(opcode_2)

        //literal
        16'd0:
        begin
          result<=$signed(literal_2);
          write_enable <= 1;
        end

        //addl
        16'd1:
        begin
          result<=operand_a + literal_2;
          write_enable <= 1;
        end

        //store
        16'd2:
        begin
        end

        //call
        16'd3:
        begin
          result <= program_counter_2 + 1;
          write_enable <= 1;
          program_counter <= literal_2;
          state <= instruction_fetch;
        end

        //stop
        16'd4:
        begin
        state <= stop;
        end

        //literal_hi
        16'd5:
        begin
          result<= {literal_2, operand_a[15:0]};
          write_enable <= 1;
        end

        //wait_clocks
        16'd6:
        begin
          timer <= operand_a;
          state <= wait_state;
        end

        //load
        16'd7:
        begin
          state <= load;
        end

        //unsigned_shift_right
        16'd8:
        begin
          if(operand_b < 32) begin
            result <= operand_a >> operand_b;
            carry <= operand_a << (32-operand_b);
          end else begin
            result <= 0;
            carry <= operand_a;
          end
          write_enable <= 1;
        end

        //unsigned_greater
        16'd9:
        begin
          result <= $unsigned(operand_a) > $unsigned(operand_b);
          write_enable <= 1;
        end

        //jmp_if_false
        16'd10:
        begin
          if (operand_a == 0) begin
            program_counter <= literal_2;
            state <= instruction_fetch;
          end
        end

        //add
        16'd11:
        begin
          long_result = operand_a + operand_b;
          result <= long_result[31:0];
          carry[0] <= long_result[32];
          write_enable <= 1;
        end

        //write
        16'd12:
        begin
          state <= write;
          write_output <= operand_a;
          write_value <= operand_b;
        end

        //goto
        16'd13:
        begin
          program_counter <= literal_2;
          state <= instruction_fetch;
        end

        //return
        16'd14:
        begin
          program_counter <= operand_a;
          state <= instruction_fetch;
        end

        //read
        16'd15:
        begin
          state <= read;
          read_input <= operand_a;
        end

        //subtract
        16'd16:
        begin
          long_result = operand_a + (~operand_b) + 1;
          result <= long_result[31:0];
          carry[0] <= ~long_result[32];
          write_enable <= 1;
        end

        //equal
        16'd17:
        begin
          result <= operand_a == operand_b;
          write_enable <= 1;
        end

      endcase

    end

    read:
    begin
      case(read_input)
      2:
      begin
        s_input_eth_in_ack <= 1;
        if (s_input_eth_in_ack && input_eth_in_stb) begin
          result <= input_eth_in;
          write_enable <= 1;
          s_input_eth_in_ack <= 0;
          state <= execute;
        end
      end
      endcase
    end

    write:
    begin
      case(write_output)
      0:
      begin
        s_output_audio_out_stb <= 1;
        s_output_audio_out <= write_value;
        if (output_audio_out_ack && s_output_audio_out_stb) begin
          s_output_audio_out_stb <= 0;
          state <= execute;
        end
      end
      1:
      begin
        s_output_eth_out_stb <= 1;
        s_output_eth_out <= write_value;
        if (output_eth_out_ack && s_output_eth_out_stb) begin
          s_output_eth_out_stb <= 0;
          state <= execute;
        end
      end
      endcase
    end

    load:
    begin
        result <= load_data;
        write_enable <= 1;
        state <= execute;
    end

    wait_state:
    begin
      if (timer) begin
        timer <= timer - 1;
      end else begin
        state <= execute;
      end
    end

    stop:
    begin
    end

    endcase

    if (rst == 1'b1) begin
      timer <= 0;
      timer_clock <= 0;
      program_counter <= 0;
      address_z_3 <= 0;
      result <= 0;
      a = 0;
      b = 0;
      z = 0;
      state <= instruction_fetch;
      s_input_eth_in_ack <= 0;
      s_output_audio_out_stb <= 0;
      s_output_eth_out_stb <= 0;
    end
  end
  assign input_eth_in_ack = s_input_eth_in_ack;
  assign output_audio_out_stb = s_output_audio_out_stb;
  assign output_audio_out = s_output_audio_out;
  assign output_eth_out_stb = s_output_eth_out_stb;
  assign output_eth_out = s_output_eth_out;

endmodule
