//name : main_0
//input : input_rs232_rx:16
//output : output_led_r:16
//output : output_led_g:16
//output : output_led_b:16
//output : output_rs232_tx:16
//source_file : /tmp/tmpn6Oyv3/inline_c_file.c

///+============================================================================+
///|                                                                            |
///|                     This file was generated by Chips                       |
///|                                                                            |
///|                                  Chips                                     |
///|                                                                            |
///|                      http://github.com/dawsonjon/Chips-2.0                 |
///|                                                                            |
///|                                                             Python powered |
///+============================================================================+
module main_0(input_rs232_rx,input_rs232_rx_stb,output_led_r_ack,output_led_g_ack,output_led_b_ack,output_rs232_tx_ack,clk,rst,output_led_r,output_led_g,output_led_b,output_rs232_tx,output_led_r_stb,output_led_g_stb,output_led_b_stb,output_rs232_tx_stb,input_rs232_rx_ack,exception);
  integer file_count;
  parameter  stop = 3'd0,
  instruction_fetch = 3'd1,
  operand_fetch = 3'd2,
  execute = 3'd3,
  load = 3'd4,
  wait_state = 3'd5,
  read = 3'd6,
  write = 3'd7;
  input [31:0] input_rs232_rx;
  input input_rs232_rx_stb;
  input output_led_r_ack;
  input output_led_g_ack;
  input output_led_b_ack;
  input output_rs232_tx_ack;
  input clk;
  input rst;
  output [31:0] output_led_r;
  output [31:0] output_led_g;
  output [31:0] output_led_b;
  output [31:0] output_rs232_tx;
  output output_led_r_stb;
  output output_led_g_stb;
  output output_led_b_stb;
  output output_rs232_tx_stb;
  output input_rs232_rx_ack;
  reg [31:0] timer;
  reg [63:0] timer_clock;
  reg [15:0] program_counter;
  reg [15:0] program_counter_1;
  reg [15:0] program_counter_2;
  reg [44:0] instruction;
  reg [4:0] opcode_2;
  reg [3:0] a;
  reg [3:0] b;
  reg [3:0] z;
  reg write_enable;
  reg [3:0] address_a_2;
  reg [3:0] address_b_2;
  reg [3:0] address_z_2;
  reg [3:0] address_z_3;
  reg [31:0] load_data;
  reg [31:0] write_output;
  reg [31:0] write_value;
  reg [31:0] read_input;
  reg [15:0] literal_2;
  reg [31:0] a_hi;
  reg [31:0] b_hi;
  reg [31:0] a_lo;
  reg [31:0] b_lo;
  reg [63:0] long_result;
  reg [31:0] result;
  reg [15:0] address;
  reg [31:0] data_out;
  reg [31:0] data_in;
  reg [31:0] carry;
  reg [31:0] s_output_led_r_stb;
  reg [31:0] s_output_led_g_stb;
  reg [31:0] s_output_led_b_stb;
  reg [31:0] s_output_rs232_tx_stb;
  reg [31:0] s_output_led_r;
  reg [31:0] s_output_led_g;
  reg [31:0] s_output_led_b;
  reg [31:0] s_output_rs232_tx;
  reg [31:0] s_input_rs232_rx_ack;
  reg [7:0] state;
  output reg exception;
  reg [28:0] instructions [1274:0];
  reg [31:0] memory [4096:0];
  reg [31:0] registers [15:0];
  wire [31:0] operand_a;
  wire [31:0] operand_b;
  wire [31:0] register_a;
  wire [31:0] register_b;
  wire [15:0] literal;
  wire [4:0] opcode;
  wire [3:0] address_a;
  wire [3:0] address_b;
  wire [3:0] address_z;
  wire [15:0] load_address;
  wire [15:0] store_address;
  wire [31:0] store_data;
  wire  store_enable;

  //////////////////////////////////////////////////////////////////////////////
  // INSTRUCTION INITIALIZATION                                                 
  //                                                                            
  // Initialise the contents of the instruction memory                          
  //
  // Intruction Set
  // ==============
  // 0 {'literal': True, 'op': 'literal'}
  // 1 {'literal': True, 'op': 'addl'}
  // 2 {'literal': False, 'op': 'store'}
  // 3 {'literal': True, 'op': 'call'}
  // 4 {'literal': False, 'op': 'stop'}
  // 5 {'literal': False, 'op': 'load'}
  // 6 {'literal': True, 'op': 'goto'}
  // 7 {'literal': False, 'op': 'return'}
  // 8 {'literal': False, 'op': 'add'}
  // 9 {'literal': True, 'op': 'jmp_if_false'}
  // 10 {'literal': False, 'op': 'write'}
  // 11 {'literal': False, 'op': 'read'}
  // 12 {'literal': False, 'op': 'equal'}
  // 13 {'literal': False, 'op': 'shift_left'}
  // 14 {'literal': False, 'op': 'greater_equal'}
  // 15 {'literal': True, 'op': 'jmp_if_true'}
  // 16 {'literal': False, 'op': 'subtract'}
  // 17 {'literal': False, 'op': 'unsigned_greater'}
  // 18 {'literal': False, 'op': 'unsigned_shift_right'}
  // Intructions
  // ===========
  
  initial
  begin
    instructions[0] = {5'd0, 4'd3, 4'd0, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 44 {'literal': 0, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 44, 'op': 'literal'}
    instructions[1] = {5'd0, 4'd4, 4'd0, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 44 {'literal': 0, 'z': 4, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 44, 'op': 'literal'}
    instructions[2] = {5'd1, 4'd3, 4'd3, 16'd145};///tmp/tmpn6Oyv3/inline_c_file.c : 44 {'a': 3, 'literal': 145, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 44, 'op': 'addl'}
    instructions[3] = {5'd0, 4'd8, 4'd0, 16'd101};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 101, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[4] = {5'd0, 4'd2, 4'd0, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 1, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[5] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'store'}
    instructions[6] = {5'd0, 4'd8, 4'd0, 16'd110};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 110, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[7] = {5'd0, 4'd2, 4'd0, 16'd2};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 2, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[8] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'store'}
    instructions[9] = {5'd0, 4'd8, 4'd0, 16'd116};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 116, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[10] = {5'd0, 4'd2, 4'd0, 16'd3};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 3, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[11] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'store'}
    instructions[12] = {5'd0, 4'd8, 4'd0, 16'd101};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 101, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[13] = {5'd0, 4'd2, 4'd0, 16'd4};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 4, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[14] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'store'}
    instructions[15] = {5'd0, 4'd8, 4'd0, 16'd114};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 114, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[16] = {5'd0, 4'd2, 4'd0, 16'd5};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 5, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[17] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'store'}
    instructions[18] = {5'd0, 4'd8, 4'd0, 16'd32};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 32, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[19] = {5'd0, 4'd2, 4'd0, 16'd6};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 6, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[20] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'store'}
    instructions[21] = {5'd0, 4'd8, 4'd0, 16'd114};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 114, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[22] = {5'd0, 4'd2, 4'd0, 16'd7};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 7, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[23] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'store'}
    instructions[24] = {5'd0, 4'd8, 4'd0, 16'd101};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 101, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[25] = {5'd0, 4'd2, 4'd0, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 8, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[26] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'store'}
    instructions[27] = {5'd0, 4'd8, 4'd0, 16'd100};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 100, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[28] = {5'd0, 4'd2, 4'd0, 16'd9};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 9, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[29] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'store'}
    instructions[30] = {5'd0, 4'd8, 4'd0, 16'd32};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 32, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[31] = {5'd0, 4'd2, 4'd0, 16'd10};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 10, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[32] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'store'}
    instructions[33] = {5'd0, 4'd8, 4'd0, 16'd108};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 108, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[34] = {5'd0, 4'd2, 4'd0, 16'd11};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 11, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[35] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'store'}
    instructions[36] = {5'd0, 4'd8, 4'd0, 16'd101};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 101, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[37] = {5'd0, 4'd2, 4'd0, 16'd12};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 12, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[38] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'store'}
    instructions[39] = {5'd0, 4'd8, 4'd0, 16'd118};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 118, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[40] = {5'd0, 4'd2, 4'd0, 16'd13};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 13, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[41] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'store'}
    instructions[42] = {5'd0, 4'd8, 4'd0, 16'd101};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 101, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[43] = {5'd0, 4'd2, 4'd0, 16'd14};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 14, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[44] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'store'}
    instructions[45] = {5'd0, 4'd8, 4'd0, 16'd108};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 108, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[46] = {5'd0, 4'd2, 4'd0, 16'd15};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 15, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[47] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'store'}
    instructions[48] = {5'd0, 4'd8, 4'd0, 16'd32};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 32, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[49] = {5'd0, 4'd2, 4'd0, 16'd16};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 16, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[50] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'store'}
    instructions[51] = {5'd0, 4'd8, 4'd0, 16'd40};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 40, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[52] = {5'd0, 4'd2, 4'd0, 16'd17};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 17, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[53] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'store'}
    instructions[54] = {5'd0, 4'd8, 4'd0, 16'd104};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 104, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[55] = {5'd0, 4'd2, 4'd0, 16'd18};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 18, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[56] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'store'}
    instructions[57] = {5'd0, 4'd8, 4'd0, 16'd101};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 101, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[58] = {5'd0, 4'd2, 4'd0, 16'd19};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 19, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[59] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'store'}
    instructions[60] = {5'd0, 4'd8, 4'd0, 16'd120};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 120, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[61] = {5'd0, 4'd2, 4'd0, 16'd20};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 20, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[62] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'store'}
    instructions[63] = {5'd0, 4'd8, 4'd0, 16'd32};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 32, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[64] = {5'd0, 4'd2, 4'd0, 16'd21};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 21, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[65] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'store'}
    instructions[66] = {5'd0, 4'd8, 4'd0, 16'd48};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 48, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[67] = {5'd0, 4'd2, 4'd0, 16'd22};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 22, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[68] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'store'}
    instructions[69] = {5'd0, 4'd8, 4'd0, 16'd45};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 45, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[70] = {5'd0, 4'd2, 4'd0, 16'd23};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 23, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[71] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'store'}
    instructions[72] = {5'd0, 4'd8, 4'd0, 16'd70};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 70, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[73] = {5'd0, 4'd2, 4'd0, 16'd24};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 24, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[74] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'store'}
    instructions[75] = {5'd0, 4'd8, 4'd0, 16'd70};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 70, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[76] = {5'd0, 4'd2, 4'd0, 16'd25};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 25, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[77] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'store'}
    instructions[78] = {5'd0, 4'd8, 4'd0, 16'd41};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 41, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[79] = {5'd0, 4'd2, 4'd0, 16'd26};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 26, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[80] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'store'}
    instructions[81] = {5'd0, 4'd8, 4'd0, 16'd10};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 10, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[82] = {5'd0, 4'd2, 4'd0, 16'd27};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 27, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[83] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'store'}
    instructions[84] = {5'd0, 4'd8, 4'd0, 16'd32};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 32, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[85] = {5'd0, 4'd2, 4'd0, 16'd28};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 28, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[86] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'store'}
    instructions[87] = {5'd0, 4'd8, 4'd0, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 0, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[88] = {5'd0, 4'd2, 4'd0, 16'd29};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 29, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[89] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'store'}
    instructions[90] = {5'd0, 4'd8, 4'd0, 16'd10};///tmp/tmpn6Oyv3/inline_c_file.c : 35 {'literal': 10, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 35, 'op': 'literal'}
    instructions[91] = {5'd0, 4'd2, 4'd0, 16'd31};///tmp/tmpn6Oyv3/inline_c_file.c : 35 {'literal': 31, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 35, 'op': 'literal'}
    instructions[92] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 35 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 35, 'op': 'store'}
    instructions[93] = {5'd0, 4'd8, 4'd0, 16'd32};///tmp/tmpn6Oyv3/inline_c_file.c : 35 {'literal': 32, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 35, 'op': 'literal'}
    instructions[94] = {5'd0, 4'd2, 4'd0, 16'd32};///tmp/tmpn6Oyv3/inline_c_file.c : 35 {'literal': 32, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 35, 'op': 'literal'}
    instructions[95] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 35 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 35, 'op': 'store'}
    instructions[96] = {5'd0, 4'd8, 4'd0, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 35 {'literal': 0, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 35, 'op': 'literal'}
    instructions[97] = {5'd0, 4'd2, 4'd0, 16'd33};///tmp/tmpn6Oyv3/inline_c_file.c : 35 {'literal': 33, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 35, 'op': 'literal'}
    instructions[98] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 35 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 35, 'op': 'store'}
    instructions[99] = {5'd0, 4'd8, 4'd0, 16'd10};///tmp/tmpn6Oyv3/inline_c_file.c : 30 {'literal': 10, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 30, 'op': 'literal'}
    instructions[100] = {5'd0, 4'd2, 4'd0, 16'd34};///tmp/tmpn6Oyv3/inline_c_file.c : 30 {'literal': 34, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 30, 'op': 'literal'}
    instructions[101] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 30 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 30, 'op': 'store'}
    instructions[102] = {5'd0, 4'd8, 4'd0, 16'd32};///tmp/tmpn6Oyv3/inline_c_file.c : 30 {'literal': 32, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 30, 'op': 'literal'}
    instructions[103] = {5'd0, 4'd2, 4'd0, 16'd35};///tmp/tmpn6Oyv3/inline_c_file.c : 30 {'literal': 35, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 30, 'op': 'literal'}
    instructions[104] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 30 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 30, 'op': 'store'}
    instructions[105] = {5'd0, 4'd8, 4'd0, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 30 {'literal': 0, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 30, 'op': 'literal'}
    instructions[106] = {5'd0, 4'd2, 4'd0, 16'd36};///tmp/tmpn6Oyv3/inline_c_file.c : 30 {'literal': 36, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 30, 'op': 'literal'}
    instructions[107] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 30 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 30, 'op': 'store'}
    instructions[108] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 4 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 4, 'op': 'literal'}
    instructions[109] = {5'd0, 4'd2, 4'd0, 16'd38};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 4 {'literal': 38, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 4, 'op': 'literal'}
    instructions[110] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 4 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 4, 'op': 'store'}
    instructions[111] = {5'd0, 4'd8, 4'd0, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 5 {'literal': 0, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 5, 'op': 'literal'}
    instructions[112] = {5'd0, 4'd2, 4'd0, 16'd39};///tmp/tmpn6Oyv3/inline_c_file.c : 5 {'literal': 39, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 5, 'op': 'literal'}
    instructions[113] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 5 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 5, 'op': 'store'}
    instructions[114] = {5'd0, 4'd8, 4'd0, 16'd101};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 101, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[115] = {5'd0, 4'd2, 4'd0, 16'd41};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 41, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[116] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'store'}
    instructions[117] = {5'd0, 4'd8, 4'd0, 16'd110};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 110, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[118] = {5'd0, 4'd2, 4'd0, 16'd42};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 42, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[119] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'store'}
    instructions[120] = {5'd0, 4'd8, 4'd0, 16'd116};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 116, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[121] = {5'd0, 4'd2, 4'd0, 16'd43};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 43, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[122] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'store'}
    instructions[123] = {5'd0, 4'd8, 4'd0, 16'd101};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 101, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[124] = {5'd0, 4'd2, 4'd0, 16'd44};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 44, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[125] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'store'}
    instructions[126] = {5'd0, 4'd8, 4'd0, 16'd114};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 114, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[127] = {5'd0, 4'd2, 4'd0, 16'd45};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 45, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[128] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'store'}
    instructions[129] = {5'd0, 4'd8, 4'd0, 16'd32};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 32, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[130] = {5'd0, 4'd2, 4'd0, 16'd46};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 46, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[131] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'store'}
    instructions[132] = {5'd0, 4'd8, 4'd0, 16'd98};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 98, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[133] = {5'd0, 4'd2, 4'd0, 16'd47};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 47, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[134] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'store'}
    instructions[135] = {5'd0, 4'd8, 4'd0, 16'd108};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 108, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[136] = {5'd0, 4'd2, 4'd0, 16'd48};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 48, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[137] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'store'}
    instructions[138] = {5'd0, 4'd8, 4'd0, 16'd117};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 117, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[139] = {5'd0, 4'd2, 4'd0, 16'd49};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 49, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[140] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'store'}
    instructions[141] = {5'd0, 4'd8, 4'd0, 16'd101};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 101, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[142] = {5'd0, 4'd2, 4'd0, 16'd50};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 50, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[143] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'store'}
    instructions[144] = {5'd0, 4'd8, 4'd0, 16'd32};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 32, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[145] = {5'd0, 4'd2, 4'd0, 16'd51};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 51, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[146] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'store'}
    instructions[147] = {5'd0, 4'd8, 4'd0, 16'd108};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 108, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[148] = {5'd0, 4'd2, 4'd0, 16'd52};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 52, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[149] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'store'}
    instructions[150] = {5'd0, 4'd8, 4'd0, 16'd101};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 101, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[151] = {5'd0, 4'd2, 4'd0, 16'd53};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 53, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[152] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'store'}
    instructions[153] = {5'd0, 4'd8, 4'd0, 16'd118};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 118, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[154] = {5'd0, 4'd2, 4'd0, 16'd54};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 54, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[155] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'store'}
    instructions[156] = {5'd0, 4'd8, 4'd0, 16'd101};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 101, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[157] = {5'd0, 4'd2, 4'd0, 16'd55};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 55, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[158] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'store'}
    instructions[159] = {5'd0, 4'd8, 4'd0, 16'd108};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 108, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[160] = {5'd0, 4'd2, 4'd0, 16'd56};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 56, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[161] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'store'}
    instructions[162] = {5'd0, 4'd8, 4'd0, 16'd32};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 32, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[163] = {5'd0, 4'd2, 4'd0, 16'd57};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 57, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[164] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'store'}
    instructions[165] = {5'd0, 4'd8, 4'd0, 16'd40};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 40, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[166] = {5'd0, 4'd2, 4'd0, 16'd58};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 58, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[167] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'store'}
    instructions[168] = {5'd0, 4'd8, 4'd0, 16'd104};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 104, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[169] = {5'd0, 4'd2, 4'd0, 16'd59};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 59, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[170] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'store'}
    instructions[171] = {5'd0, 4'd8, 4'd0, 16'd101};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 101, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[172] = {5'd0, 4'd2, 4'd0, 16'd60};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 60, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[173] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'store'}
    instructions[174] = {5'd0, 4'd8, 4'd0, 16'd120};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 120, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[175] = {5'd0, 4'd2, 4'd0, 16'd61};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 61, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[176] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'store'}
    instructions[177] = {5'd0, 4'd8, 4'd0, 16'd32};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 32, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[178] = {5'd0, 4'd2, 4'd0, 16'd62};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 62, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[179] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'store'}
    instructions[180] = {5'd0, 4'd8, 4'd0, 16'd48};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 48, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[181] = {5'd0, 4'd2, 4'd0, 16'd63};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 63, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[182] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'store'}
    instructions[183] = {5'd0, 4'd8, 4'd0, 16'd45};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 45, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[184] = {5'd0, 4'd2, 4'd0, 16'd64};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 64, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[185] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'store'}
    instructions[186] = {5'd0, 4'd8, 4'd0, 16'd70};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 70, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[187] = {5'd0, 4'd2, 4'd0, 16'd65};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 65, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[188] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'store'}
    instructions[189] = {5'd0, 4'd8, 4'd0, 16'd70};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 70, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[190] = {5'd0, 4'd2, 4'd0, 16'd66};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 66, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[191] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'store'}
    instructions[192] = {5'd0, 4'd8, 4'd0, 16'd41};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 41, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[193] = {5'd0, 4'd2, 4'd0, 16'd67};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 67, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[194] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'store'}
    instructions[195] = {5'd0, 4'd8, 4'd0, 16'd10};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 10, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[196] = {5'd0, 4'd2, 4'd0, 16'd68};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 68, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[197] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'store'}
    instructions[198] = {5'd0, 4'd8, 4'd0, 16'd32};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 32, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[199] = {5'd0, 4'd2, 4'd0, 16'd69};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 69, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[200] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'store'}
    instructions[201] = {5'd0, 4'd8, 4'd0, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 0, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[202] = {5'd0, 4'd2, 4'd0, 16'd70};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 70, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[203] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'store'}
    instructions[204] = {5'd0, 4'd8, 4'd0, 16'd67};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 67, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[205] = {5'd0, 4'd2, 4'd0, 16'd71};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 71, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[206] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'store'}
    instructions[207] = {5'd0, 4'd8, 4'd0, 16'd104};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 104, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[208] = {5'd0, 4'd2, 4'd0, 16'd72};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 72, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[209] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'store'}
    instructions[210] = {5'd0, 4'd8, 4'd0, 16'd105};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 105, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[211] = {5'd0, 4'd2, 4'd0, 16'd73};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 73, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[212] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'store'}
    instructions[213] = {5'd0, 4'd8, 4'd0, 16'd112};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 112, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[214] = {5'd0, 4'd2, 4'd0, 16'd74};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 74, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[215] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'store'}
    instructions[216] = {5'd0, 4'd8, 4'd0, 16'd115};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 115, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[217] = {5'd0, 4'd2, 4'd0, 16'd75};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 75, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[218] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'store'}
    instructions[219] = {5'd0, 4'd8, 4'd0, 16'd32};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 32, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[220] = {5'd0, 4'd2, 4'd0, 16'd76};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 76, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[221] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'store'}
    instructions[222] = {5'd0, 4'd8, 4'd0, 16'd68};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 68, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[223] = {5'd0, 4'd2, 4'd0, 16'd77};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 77, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[224] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'store'}
    instructions[225] = {5'd0, 4'd8, 4'd0, 16'd101};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 101, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[226] = {5'd0, 4'd2, 4'd0, 16'd78};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 78, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[227] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'store'}
    instructions[228] = {5'd0, 4'd8, 4'd0, 16'd109};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 109, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[229] = {5'd0, 4'd2, 4'd0, 16'd79};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 79, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[230] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'store'}
    instructions[231] = {5'd0, 4'd8, 4'd0, 16'd111};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 111, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[232] = {5'd0, 4'd2, 4'd0, 16'd80};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 80, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[233] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'store'}
    instructions[234] = {5'd0, 4'd8, 4'd0, 16'd32};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 32, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[235] = {5'd0, 4'd2, 4'd0, 16'd81};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 81, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[236] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'store'}
    instructions[237] = {5'd0, 4'd8, 4'd0, 16'd116};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 116, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[238] = {5'd0, 4'd2, 4'd0, 16'd82};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 82, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[239] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'store'}
    instructions[240] = {5'd0, 4'd8, 4'd0, 16'd114};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 114, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[241] = {5'd0, 4'd2, 4'd0, 16'd83};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 83, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[242] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'store'}
    instructions[243] = {5'd0, 4'd8, 4'd0, 16'd105};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 105, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[244] = {5'd0, 4'd2, 4'd0, 16'd84};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 84, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[245] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'store'}
    instructions[246] = {5'd0, 4'd8, 4'd0, 16'd45};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 45, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[247] = {5'd0, 4'd2, 4'd0, 16'd85};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 85, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[248] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'store'}
    instructions[249] = {5'd0, 4'd8, 4'd0, 16'd99};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 99, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[250] = {5'd0, 4'd2, 4'd0, 16'd86};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 86, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[251] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'store'}
    instructions[252] = {5'd0, 4'd8, 4'd0, 16'd111};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 111, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[253] = {5'd0, 4'd2, 4'd0, 16'd87};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 87, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[254] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'store'}
    instructions[255] = {5'd0, 4'd8, 4'd0, 16'd108};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 108, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[256] = {5'd0, 4'd2, 4'd0, 16'd88};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 88, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[257] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'store'}
    instructions[258] = {5'd0, 4'd8, 4'd0, 16'd111};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 111, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[259] = {5'd0, 4'd2, 4'd0, 16'd89};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 89, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[260] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'store'}
    instructions[261] = {5'd0, 4'd8, 4'd0, 16'd114};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 114, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[262] = {5'd0, 4'd2, 4'd0, 16'd90};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 90, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[263] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'store'}
    instructions[264] = {5'd0, 4'd8, 4'd0, 16'd32};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 32, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[265] = {5'd0, 4'd2, 4'd0, 16'd91};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 91, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[266] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'store'}
    instructions[267] = {5'd0, 4'd8, 4'd0, 16'd76};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 76, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[268] = {5'd0, 4'd2, 4'd0, 16'd92};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 92, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[269] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'store'}
    instructions[270] = {5'd0, 4'd8, 4'd0, 16'd69};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 69, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[271] = {5'd0, 4'd2, 4'd0, 16'd93};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 93, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[272] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'store'}
    instructions[273] = {5'd0, 4'd8, 4'd0, 16'd68};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 68, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[274] = {5'd0, 4'd2, 4'd0, 16'd94};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 94, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[275] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'store'}
    instructions[276] = {5'd0, 4'd8, 4'd0, 16'd32};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 32, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[277] = {5'd0, 4'd2, 4'd0, 16'd95};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 95, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[278] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'store'}
    instructions[279] = {5'd0, 4'd8, 4'd0, 16'd101};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 101, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[280] = {5'd0, 4'd2, 4'd0, 16'd96};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 96, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[281] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'store'}
    instructions[282] = {5'd0, 4'd8, 4'd0, 16'd120};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 120, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[283] = {5'd0, 4'd2, 4'd0, 16'd97};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 97, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[284] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'store'}
    instructions[285] = {5'd0, 4'd8, 4'd0, 16'd97};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 97, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[286] = {5'd0, 4'd2, 4'd0, 16'd98};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 98, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[287] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'store'}
    instructions[288] = {5'd0, 4'd8, 4'd0, 16'd109};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 109, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[289] = {5'd0, 4'd2, 4'd0, 16'd99};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 99, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[290] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'store'}
    instructions[291] = {5'd0, 4'd8, 4'd0, 16'd112};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 112, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[292] = {5'd0, 4'd2, 4'd0, 16'd100};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 100, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[293] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'store'}
    instructions[294] = {5'd0, 4'd8, 4'd0, 16'd108};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 108, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[295] = {5'd0, 4'd2, 4'd0, 16'd101};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 101, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[296] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'store'}
    instructions[297] = {5'd0, 4'd8, 4'd0, 16'd101};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 101, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[298] = {5'd0, 4'd2, 4'd0, 16'd102};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 102, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[299] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'store'}
    instructions[300] = {5'd0, 4'd8, 4'd0, 16'd10};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 10, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[301] = {5'd0, 4'd2, 4'd0, 16'd103};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 103, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[302] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'store'}
    instructions[303] = {5'd0, 4'd8, 4'd0, 16'd32};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 32, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[304] = {5'd0, 4'd2, 4'd0, 16'd104};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 104, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[305] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'store'}
    instructions[306] = {5'd0, 4'd8, 4'd0, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 0, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[307] = {5'd0, 4'd2, 4'd0, 16'd105};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 105, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[308] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'store'}
    instructions[309] = {5'd0, 4'd8, 4'd0, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 6 {'literal': 1, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 6, 'op': 'literal'}
    instructions[310] = {5'd0, 4'd2, 4'd0, 16'd106};///tmp/tmpn6Oyv3/inline_c_file.c : 6 {'literal': 106, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 6, 'op': 'literal'}
    instructions[311] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 6 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 6, 'op': 'store'}
    instructions[312] = {5'd0, 4'd8, 4'd0, 16'd2};///tmp/tmpn6Oyv3/inline_c_file.c : 7 {'literal': 2, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 7, 'op': 'literal'}
    instructions[313] = {5'd0, 4'd2, 4'd0, 16'd107};///tmp/tmpn6Oyv3/inline_c_file.c : 7 {'literal': 107, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 7, 'op': 'literal'}
    instructions[314] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 7 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 7, 'op': 'store'}
    instructions[315] = {5'd0, 4'd8, 4'd0, 16'd10};///tmp/tmpn6Oyv3/inline_c_file.c : 40 {'literal': 10, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 40, 'op': 'literal'}
    instructions[316] = {5'd0, 4'd2, 4'd0, 16'd108};///tmp/tmpn6Oyv3/inline_c_file.c : 40 {'literal': 108, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 40, 'op': 'literal'}
    instructions[317] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 40 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 40, 'op': 'store'}
    instructions[318] = {5'd0, 4'd8, 4'd0, 16'd32};///tmp/tmpn6Oyv3/inline_c_file.c : 40 {'literal': 32, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 40, 'op': 'literal'}
    instructions[319] = {5'd0, 4'd2, 4'd0, 16'd109};///tmp/tmpn6Oyv3/inline_c_file.c : 40 {'literal': 109, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 40, 'op': 'literal'}
    instructions[320] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 40 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 40, 'op': 'store'}
    instructions[321] = {5'd0, 4'd8, 4'd0, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 40 {'literal': 0, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 40, 'op': 'literal'}
    instructions[322] = {5'd0, 4'd2, 4'd0, 16'd110};///tmp/tmpn6Oyv3/inline_c_file.c : 40 {'literal': 110, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 40, 'op': 'literal'}
    instructions[323] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 40 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 40, 'op': 'store'}
    instructions[324] = {5'd0, 4'd8, 4'd0, 16'd3};///tmp/tmpn6Oyv3/inline_c_file.c : 8 {'literal': 3, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 8, 'op': 'literal'}
    instructions[325] = {5'd0, 4'd2, 4'd0, 16'd111};///tmp/tmpn6Oyv3/inline_c_file.c : 8 {'literal': 111, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 8, 'op': 'literal'}
    instructions[326] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 8 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 8, 'op': 'store'}
    instructions[327] = {5'd0, 4'd8, 4'd0, 16'd4};///tmp/tmpn6Oyv3/inline_c_file.c : 9 {'literal': 4, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 9, 'op': 'literal'}
    instructions[328] = {5'd0, 4'd2, 4'd0, 16'd112};///tmp/tmpn6Oyv3/inline_c_file.c : 9 {'literal': 112, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 9, 'op': 'literal'}
    instructions[329] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 9 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 9, 'op': 'store'}
    instructions[330] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 5 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 5, 'op': 'literal'}
    instructions[331] = {5'd0, 4'd2, 4'd0, 16'd113};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 5 {'literal': 113, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 5, 'op': 'literal'}
    instructions[332] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 5 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 5, 'op': 'store'}
    instructions[333] = {5'd0, 4'd8, 4'd0, 16'd101};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 101, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[334] = {5'd0, 4'd2, 4'd0, 16'd114};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 114, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[335] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'store'}
    instructions[336] = {5'd0, 4'd8, 4'd0, 16'd110};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 110, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[337] = {5'd0, 4'd2, 4'd0, 16'd115};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 115, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[338] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'store'}
    instructions[339] = {5'd0, 4'd8, 4'd0, 16'd116};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 116, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[340] = {5'd0, 4'd2, 4'd0, 16'd116};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 116, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[341] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'store'}
    instructions[342] = {5'd0, 4'd8, 4'd0, 16'd101};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 101, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[343] = {5'd0, 4'd2, 4'd0, 16'd117};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 117, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[344] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'store'}
    instructions[345] = {5'd0, 4'd8, 4'd0, 16'd114};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 114, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[346] = {5'd0, 4'd2, 4'd0, 16'd118};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 118, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[347] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'store'}
    instructions[348] = {5'd0, 4'd8, 4'd0, 16'd32};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 32, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[349] = {5'd0, 4'd2, 4'd0, 16'd119};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 119, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[350] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'store'}
    instructions[351] = {5'd0, 4'd8, 4'd0, 16'd103};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 103, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[352] = {5'd0, 4'd2, 4'd0, 16'd120};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 120, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[353] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'store'}
    instructions[354] = {5'd0, 4'd8, 4'd0, 16'd114};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 114, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[355] = {5'd0, 4'd2, 4'd0, 16'd121};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 121, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[356] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'store'}
    instructions[357] = {5'd0, 4'd8, 4'd0, 16'd101};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 101, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[358] = {5'd0, 4'd2, 4'd0, 16'd122};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 122, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[359] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'store'}
    instructions[360] = {5'd0, 4'd8, 4'd0, 16'd101};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 101, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[361] = {5'd0, 4'd2, 4'd0, 16'd123};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 123, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[362] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'store'}
    instructions[363] = {5'd0, 4'd8, 4'd0, 16'd110};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 110, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[364] = {5'd0, 4'd2, 4'd0, 16'd124};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 124, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[365] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'store'}
    instructions[366] = {5'd0, 4'd8, 4'd0, 16'd32};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 32, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[367] = {5'd0, 4'd2, 4'd0, 16'd125};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 125, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[368] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'store'}
    instructions[369] = {5'd0, 4'd8, 4'd0, 16'd108};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 108, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[370] = {5'd0, 4'd2, 4'd0, 16'd126};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 126, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[371] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'store'}
    instructions[372] = {5'd0, 4'd8, 4'd0, 16'd101};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 101, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[373] = {5'd0, 4'd2, 4'd0, 16'd127};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 127, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[374] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'store'}
    instructions[375] = {5'd0, 4'd8, 4'd0, 16'd118};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 118, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[376] = {5'd0, 4'd2, 4'd0, 16'd128};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 128, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[377] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'store'}
    instructions[378] = {5'd0, 4'd8, 4'd0, 16'd101};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 101, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[379] = {5'd0, 4'd2, 4'd0, 16'd129};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 129, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[380] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'store'}
    instructions[381] = {5'd0, 4'd8, 4'd0, 16'd108};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 108, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[382] = {5'd0, 4'd2, 4'd0, 16'd130};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 130, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[383] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'store'}
    instructions[384] = {5'd0, 4'd8, 4'd0, 16'd32};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 32, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[385] = {5'd0, 4'd2, 4'd0, 16'd131};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 131, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[386] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'store'}
    instructions[387] = {5'd0, 4'd8, 4'd0, 16'd40};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 40, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[388] = {5'd0, 4'd2, 4'd0, 16'd132};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 132, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[389] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'store'}
    instructions[390] = {5'd0, 4'd8, 4'd0, 16'd104};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 104, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[391] = {5'd0, 4'd2, 4'd0, 16'd133};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 133, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[392] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'store'}
    instructions[393] = {5'd0, 4'd8, 4'd0, 16'd101};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 101, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[394] = {5'd0, 4'd2, 4'd0, 16'd134};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 134, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[395] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'store'}
    instructions[396] = {5'd0, 4'd8, 4'd0, 16'd120};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 120, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[397] = {5'd0, 4'd2, 4'd0, 16'd135};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 135, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[398] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'store'}
    instructions[399] = {5'd0, 4'd8, 4'd0, 16'd32};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 32, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[400] = {5'd0, 4'd2, 4'd0, 16'd136};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 136, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[401] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'store'}
    instructions[402] = {5'd0, 4'd8, 4'd0, 16'd48};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 48, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[403] = {5'd0, 4'd2, 4'd0, 16'd137};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 137, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[404] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'store'}
    instructions[405] = {5'd0, 4'd8, 4'd0, 16'd45};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 45, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[406] = {5'd0, 4'd2, 4'd0, 16'd138};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 138, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[407] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'store'}
    instructions[408] = {5'd0, 4'd8, 4'd0, 16'd70};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 70, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[409] = {5'd0, 4'd2, 4'd0, 16'd139};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 139, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[410] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'store'}
    instructions[411] = {5'd0, 4'd8, 4'd0, 16'd70};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 70, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[412] = {5'd0, 4'd2, 4'd0, 16'd140};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 140, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[413] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'store'}
    instructions[414] = {5'd0, 4'd8, 4'd0, 16'd41};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 41, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[415] = {5'd0, 4'd2, 4'd0, 16'd141};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 141, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[416] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'store'}
    instructions[417] = {5'd0, 4'd8, 4'd0, 16'd10};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 10, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[418] = {5'd0, 4'd2, 4'd0, 16'd142};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 142, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[419] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'store'}
    instructions[420] = {5'd0, 4'd8, 4'd0, 16'd32};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 32, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[421] = {5'd0, 4'd2, 4'd0, 16'd143};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 143, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[422] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'store'}
    instructions[423] = {5'd0, 4'd8, 4'd0, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 0, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[424] = {5'd0, 4'd2, 4'd0, 16'd144};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 144, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[425] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'store'}
    instructions[426] = {5'd1, 4'd7, 4'd4, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 44 {'a': 4, 'literal': 0, 'z': 7, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 44, 'op': 'addl'}
    instructions[427] = {5'd1, 4'd4, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 44 {'a': 3, 'literal': 0, 'z': 4, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 44, 'op': 'addl'}
    instructions[428] = {5'd3, 4'd6, 4'd0, 16'd430};///tmp/tmpn6Oyv3/inline_c_file.c : 44 {'z': 6, 'label': 430, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 44, 'op': 'call'}
    instructions[429] = {5'd4, 4'd0, 4'd0, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 44 {'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 44, 'op': 'stop'}
    instructions[430] = {5'd1, 4'd3, 4'd3, 16'd137};///tmp/tmpn6Oyv3/inline_c_file.c : 17 {'a': 3, 'literal': 137, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 17, 'op': 'addl'}
    instructions[431] = {5'd0, 4'd8, 4'd0, 16'd111};///tmp/tmpn6Oyv3/inline_c_file.c : 18 {'literal': 111, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 18, 'op': 'literal'}
    instructions[432] = {5'd1, 4'd2, 4'd8, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 18 {'a': 8, 'literal': 0, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 18, 'op': 'addl'}
    instructions[433] = {5'd5, 4'd8, 4'd2, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 18 {'a': 2, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 18, 'op': 'load'}
    instructions[434] = {5'd0, 4'd2, 4'd0, 16'd113};///tmp/tmpn6Oyv3/inline_c_file.c : 18 {'literal': 113, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 18, 'op': 'literal'}
    instructions[435] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 18 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 18, 'op': 'store'}
    instructions[436] = {5'd0, 4'd8, 4'd0, 16'd112};///tmp/tmpn6Oyv3/inline_c_file.c : 19 {'literal': 112, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 19, 'op': 'literal'}
    instructions[437] = {5'd1, 4'd2, 4'd8, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 19 {'a': 8, 'literal': 0, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 19, 'op': 'addl'}
    instructions[438] = {5'd5, 4'd8, 4'd2, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 19 {'a': 2, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 19, 'op': 'load'}
    instructions[439] = {5'd0, 4'd2, 4'd0, 16'd38};///tmp/tmpn6Oyv3/inline_c_file.c : 19 {'literal': 38, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 19, 'op': 'literal'}
    instructions[440] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 19 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 19, 'op': 'store'}
    instructions[441] = {5'd2, 4'd0, 4'd3, 16'd6};///tmp/tmpn6Oyv3/inline_c_file.c : 23 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 23, 'op': 'store'}
    instructions[442] = {5'd1, 4'd3, 4'd3, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 23 {'a': 3, 'literal': 1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 23, 'op': 'addl'}
    instructions[443] = {5'd2, 4'd0, 4'd3, 16'd7};///tmp/tmpn6Oyv3/inline_c_file.c : 23 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 23, 'op': 'store'}
    instructions[444] = {5'd1, 4'd3, 4'd3, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 23 {'a': 3, 'literal': 1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 23, 'op': 'addl'}
    instructions[445] = {5'd0, 4'd8, 4'd0, 16'd71};///tmp/tmpn6Oyv3/inline_c_file.c : 24 {'literal': 71, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 24, 'op': 'literal'}
    instructions[446] = {5'd2, 4'd0, 4'd3, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 23 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 23, 'op': 'store'}
    instructions[447] = {5'd1, 4'd3, 4'd3, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 23 {'a': 3, 'literal': 1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 23, 'op': 'addl'}
    instructions[448] = {5'd1, 4'd7, 4'd4, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 23 {'a': 4, 'literal': 0, 'z': 7, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 23, 'op': 'addl'}
    instructions[449] = {5'd1, 4'd4, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 23 {'a': 3, 'literal': 0, 'z': 4, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 23, 'op': 'addl'}
    instructions[450] = {5'd3, 4'd6, 4'd0, 16'd687};///tmp/tmpn6Oyv3/inline_c_file.c : 23 {'z': 6, 'label': 687, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 23, 'op': 'call'}
    instructions[451] = {5'd1, 4'd3, 4'd3, -16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 23 {'a': 3, 'literal': -1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 23, 'op': 'addl'}
    instructions[452] = {5'd1, 4'd3, 4'd3, -16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 23 {'a': 3, 'comment': 'pop', 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 23, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[453] = {5'd5, 4'd7, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 23 {'a': 3, 'z': 7, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 23, 'op': 'load'}
    instructions[454] = {5'd1, 4'd3, 4'd3, -16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 23 {'a': 3, 'comment': 'pop', 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 23, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[455] = {5'd5, 4'd6, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 23 {'a': 3, 'z': 6, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 23, 'op': 'load'}
    instructions[456] = {5'd1, 4'd3, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 23 {'a': 3, 'literal': 0, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 23, 'op': 'addl'}
    instructions[457] = {5'd2, 4'd0, 4'd3, 16'd6};///tmp/tmpn6Oyv3/inline_c_file.c : 26 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 26, 'op': 'store'}
    instructions[458] = {5'd1, 4'd3, 4'd3, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 26 {'a': 3, 'literal': 1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 26, 'op': 'addl'}
    instructions[459] = {5'd2, 4'd0, 4'd3, 16'd7};///tmp/tmpn6Oyv3/inline_c_file.c : 26 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 26, 'op': 'store'}
    instructions[460] = {5'd1, 4'd3, 4'd3, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 26 {'a': 3, 'literal': 1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 26, 'op': 'addl'}
    instructions[461] = {5'd0, 4'd8, 4'd0, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 27 {'literal': 1, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 27, 'op': 'literal'}
    instructions[462] = {5'd2, 4'd0, 4'd3, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 26 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 26, 'op': 'store'}
    instructions[463] = {5'd1, 4'd3, 4'd3, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 26 {'a': 3, 'literal': 1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 26, 'op': 'addl'}
    instructions[464] = {5'd1, 4'd7, 4'd4, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 26 {'a': 4, 'literal': 0, 'z': 7, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 26, 'op': 'addl'}
    instructions[465] = {5'd1, 4'd4, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 26 {'a': 3, 'literal': 0, 'z': 4, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 26, 'op': 'addl'}
    instructions[466] = {5'd3, 4'd6, 4'd0, 16'd687};///tmp/tmpn6Oyv3/inline_c_file.c : 26 {'z': 6, 'label': 687, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 26, 'op': 'call'}
    instructions[467] = {5'd1, 4'd3, 4'd3, -16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 26 {'a': 3, 'literal': -1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 26, 'op': 'addl'}
    instructions[468] = {5'd1, 4'd3, 4'd3, -16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 26 {'a': 3, 'comment': 'pop', 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 26, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[469] = {5'd5, 4'd7, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 26 {'a': 3, 'z': 7, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 26, 'op': 'load'}
    instructions[470] = {5'd1, 4'd3, 4'd3, -16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 26 {'a': 3, 'comment': 'pop', 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 26, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[471] = {5'd5, 4'd6, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 26 {'a': 3, 'z': 6, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 26, 'op': 'load'}
    instructions[472] = {5'd1, 4'd3, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 26 {'a': 3, 'literal': 0, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 26, 'op': 'addl'}
    instructions[473] = {5'd2, 4'd0, 4'd3, 16'd6};///tmp/tmpn6Oyv3/inline_c_file.c : 28 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 28, 'op': 'store'}
    instructions[474] = {5'd1, 4'd3, 4'd3, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 28 {'a': 3, 'literal': 1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 28, 'op': 'addl'}
    instructions[475] = {5'd2, 4'd0, 4'd3, 16'd7};///tmp/tmpn6Oyv3/inline_c_file.c : 28 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 28, 'op': 'store'}
    instructions[476] = {5'd1, 4'd3, 4'd3, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 28 {'a': 3, 'literal': 1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 28, 'op': 'addl'}
    instructions[477] = {5'd1, 4'd7, 4'd4, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 28 {'a': 4, 'literal': 0, 'z': 7, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 28, 'op': 'addl'}
    instructions[478] = {5'd1, 4'd4, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 28 {'a': 3, 'literal': 0, 'z': 4, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 28, 'op': 'addl'}
    instructions[479] = {5'd3, 4'd6, 4'd0, 16'd778};///tmp/tmpn6Oyv3/inline_c_file.c : 28 {'z': 6, 'label': 778, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 28, 'op': 'call'}
    instructions[480] = {5'd1, 4'd3, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 28 {'a': 3, 'literal': 0, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 28, 'op': 'addl'}
    instructions[481] = {5'd1, 4'd3, 4'd3, -16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 28 {'a': 3, 'comment': 'pop', 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 28, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[482] = {5'd5, 4'd7, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 28 {'a': 3, 'z': 7, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 28, 'op': 'load'}
    instructions[483] = {5'd1, 4'd3, 4'd3, -16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 28 {'a': 3, 'comment': 'pop', 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 28, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[484] = {5'd5, 4'd6, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 28 {'a': 3, 'z': 6, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 28, 'op': 'load'}
    instructions[485] = {5'd0, 4'd2, 4'd0, 16'd37};///tmp/tmpn6Oyv3/inline_c_file.c : 28 {'literal': 37, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 28, 'op': 'literal'}
    instructions[486] = {5'd5, 4'd8, 4'd2, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 28 {'a': 2, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 28, 'op': 'load'}
    instructions[487] = {5'd1, 4'd2, 4'd4, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 28 {'a': 4, 'literal': 0, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 28, 'op': 'addl'}
    instructions[488] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 28 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 28, 'op': 'store'}
    instructions[489] = {5'd2, 4'd0, 4'd3, 16'd6};///tmp/tmpn6Oyv3/inline_c_file.c : 29 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 29, 'op': 'store'}
    instructions[490] = {5'd1, 4'd3, 4'd3, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 29 {'a': 3, 'literal': 1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 29, 'op': 'addl'}
    instructions[491] = {5'd2, 4'd0, 4'd3, 16'd7};///tmp/tmpn6Oyv3/inline_c_file.c : 29 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 29, 'op': 'store'}
    instructions[492] = {5'd1, 4'd3, 4'd3, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 29 {'a': 3, 'literal': 1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 29, 'op': 'addl'}
    instructions[493] = {5'd1, 4'd8, 4'd4, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 29 {'a': 4, 'literal': 0, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 29, 'op': 'addl'}
    instructions[494] = {5'd1, 4'd2, 4'd8, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 29 {'a': 8, 'literal': 0, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 29, 'op': 'addl'}
    instructions[495] = {5'd5, 4'd8, 4'd2, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 29 {'a': 2, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 29, 'op': 'load'}
    instructions[496] = {5'd2, 4'd0, 4'd3, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 29 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 29, 'op': 'store'}
    instructions[497] = {5'd1, 4'd3, 4'd3, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 29 {'a': 3, 'literal': 1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 29, 'op': 'addl'}
    instructions[498] = {5'd1, 4'd7, 4'd4, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 29 {'a': 4, 'literal': 0, 'z': 7, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 29, 'op': 'addl'}
    instructions[499] = {5'd1, 4'd4, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 29 {'a': 3, 'literal': 0, 'z': 4, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 29, 'op': 'addl'}
    instructions[500] = {5'd3, 4'd6, 4'd0, 16'd1079};///tmp/tmpn6Oyv3/inline_c_file.c : 29 {'z': 6, 'label': 1079, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 29, 'op': 'call'}
    instructions[501] = {5'd1, 4'd3, 4'd3, -16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 29 {'a': 3, 'literal': -1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 29, 'op': 'addl'}
    instructions[502] = {5'd1, 4'd3, 4'd3, -16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 29 {'a': 3, 'comment': 'pop', 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 29, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[503] = {5'd5, 4'd7, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 29 {'a': 3, 'z': 7, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 29, 'op': 'load'}
    instructions[504] = {5'd1, 4'd3, 4'd3, -16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 29 {'a': 3, 'comment': 'pop', 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 29, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[505] = {5'd5, 4'd6, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 29 {'a': 3, 'z': 6, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 29, 'op': 'load'}
    instructions[506] = {5'd1, 4'd3, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 29 {'a': 3, 'literal': 0, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 29, 'op': 'addl'}
    instructions[507] = {5'd2, 4'd0, 4'd3, 16'd6};///tmp/tmpn6Oyv3/inline_c_file.c : 29 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 29, 'op': 'store'}
    instructions[508] = {5'd1, 4'd3, 4'd3, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 29 {'a': 3, 'literal': 1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 29, 'op': 'addl'}
    instructions[509] = {5'd2, 4'd0, 4'd3, 16'd7};///tmp/tmpn6Oyv3/inline_c_file.c : 29 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 29, 'op': 'store'}
    instructions[510] = {5'd1, 4'd3, 4'd3, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 29 {'a': 3, 'literal': 1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 29, 'op': 'addl'}
    instructions[511] = {5'd0, 4'd8, 4'd0, 16'd34};///tmp/tmpn6Oyv3/inline_c_file.c : 30 {'literal': 34, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 30, 'op': 'literal'}
    instructions[512] = {5'd2, 4'd0, 4'd3, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 29 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 29, 'op': 'store'}
    instructions[513] = {5'd1, 4'd3, 4'd3, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 29 {'a': 3, 'literal': 1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 29, 'op': 'addl'}
    instructions[514] = {5'd1, 4'd7, 4'd4, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 29 {'a': 4, 'literal': 0, 'z': 7, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 29, 'op': 'addl'}
    instructions[515] = {5'd1, 4'd4, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 29 {'a': 3, 'literal': 0, 'z': 4, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 29, 'op': 'addl'}
    instructions[516] = {5'd3, 4'd6, 4'd0, 16'd687};///tmp/tmpn6Oyv3/inline_c_file.c : 29 {'z': 6, 'label': 687, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 29, 'op': 'call'}
    instructions[517] = {5'd1, 4'd3, 4'd3, -16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 29 {'a': 3, 'literal': -1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 29, 'op': 'addl'}
    instructions[518] = {5'd1, 4'd3, 4'd3, -16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 29 {'a': 3, 'comment': 'pop', 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 29, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[519] = {5'd5, 4'd7, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 29 {'a': 3, 'z': 7, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 29, 'op': 'load'}
    instructions[520] = {5'd1, 4'd3, 4'd3, -16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 29 {'a': 3, 'comment': 'pop', 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 29, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[521] = {5'd5, 4'd6, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 29 {'a': 3, 'z': 6, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 29, 'op': 'load'}
    instructions[522] = {5'd1, 4'd3, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 29 {'a': 3, 'literal': 0, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 29, 'op': 'addl'}
    instructions[523] = {5'd2, 4'd0, 4'd3, 16'd6};///tmp/tmpn6Oyv3/inline_c_file.c : 31 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 31, 'op': 'store'}
    instructions[524] = {5'd1, 4'd3, 4'd3, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 31 {'a': 3, 'literal': 1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 31, 'op': 'addl'}
    instructions[525] = {5'd2, 4'd0, 4'd3, 16'd7};///tmp/tmpn6Oyv3/inline_c_file.c : 31 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 31, 'op': 'store'}
    instructions[526] = {5'd1, 4'd3, 4'd3, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 31 {'a': 3, 'literal': 1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 31, 'op': 'addl'}
    instructions[527] = {5'd0, 4'd8, 4'd0, 16'd114};///tmp/tmpn6Oyv3/inline_c_file.c : 32 {'literal': 114, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 32, 'op': 'literal'}
    instructions[528] = {5'd2, 4'd0, 4'd3, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 31 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 31, 'op': 'store'}
    instructions[529] = {5'd1, 4'd3, 4'd3, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 31 {'a': 3, 'literal': 1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 31, 'op': 'addl'}
    instructions[530] = {5'd1, 4'd7, 4'd4, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 31 {'a': 4, 'literal': 0, 'z': 7, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 31, 'op': 'addl'}
    instructions[531] = {5'd1, 4'd4, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 31 {'a': 3, 'literal': 0, 'z': 4, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 31, 'op': 'addl'}
    instructions[532] = {5'd3, 4'd6, 4'd0, 16'd687};///tmp/tmpn6Oyv3/inline_c_file.c : 31 {'z': 6, 'label': 687, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 31, 'op': 'call'}
    instructions[533] = {5'd1, 4'd3, 4'd3, -16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 31 {'a': 3, 'literal': -1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 31, 'op': 'addl'}
    instructions[534] = {5'd1, 4'd3, 4'd3, -16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 31 {'a': 3, 'comment': 'pop', 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 31, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[535] = {5'd5, 4'd7, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 31 {'a': 3, 'z': 7, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 31, 'op': 'load'}
    instructions[536] = {5'd1, 4'd3, 4'd3, -16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 31 {'a': 3, 'comment': 'pop', 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 31, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[537] = {5'd5, 4'd6, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 31 {'a': 3, 'z': 6, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 31, 'op': 'load'}
    instructions[538] = {5'd1, 4'd3, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 31 {'a': 3, 'literal': 0, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 31, 'op': 'addl'}
    instructions[539] = {5'd2, 4'd0, 4'd3, 16'd6};///tmp/tmpn6Oyv3/inline_c_file.c : 33 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 33, 'op': 'store'}
    instructions[540] = {5'd1, 4'd3, 4'd3, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 33 {'a': 3, 'literal': 1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 33, 'op': 'addl'}
    instructions[541] = {5'd2, 4'd0, 4'd3, 16'd7};///tmp/tmpn6Oyv3/inline_c_file.c : 33 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 33, 'op': 'store'}
    instructions[542] = {5'd1, 4'd3, 4'd3, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 33 {'a': 3, 'literal': 1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 33, 'op': 'addl'}
    instructions[543] = {5'd1, 4'd7, 4'd4, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 33 {'a': 4, 'literal': 0, 'z': 7, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 33, 'op': 'addl'}
    instructions[544] = {5'd1, 4'd4, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 33 {'a': 3, 'literal': 0, 'z': 4, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 33, 'op': 'addl'}
    instructions[545] = {5'd3, 4'd6, 4'd0, 16'd778};///tmp/tmpn6Oyv3/inline_c_file.c : 33 {'z': 6, 'label': 778, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 33, 'op': 'call'}
    instructions[546] = {5'd1, 4'd3, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 33 {'a': 3, 'literal': 0, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 33, 'op': 'addl'}
    instructions[547] = {5'd1, 4'd3, 4'd3, -16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 33 {'a': 3, 'comment': 'pop', 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 33, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[548] = {5'd5, 4'd7, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 33 {'a': 3, 'z': 7, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 33, 'op': 'load'}
    instructions[549] = {5'd1, 4'd3, 4'd3, -16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 33 {'a': 3, 'comment': 'pop', 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 33, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[550] = {5'd5, 4'd6, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 33 {'a': 3, 'z': 6, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 33, 'op': 'load'}
    instructions[551] = {5'd0, 4'd2, 4'd0, 16'd37};///tmp/tmpn6Oyv3/inline_c_file.c : 33 {'literal': 37, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 33, 'op': 'literal'}
    instructions[552] = {5'd5, 4'd8, 4'd2, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 33 {'a': 2, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 33, 'op': 'load'}
    instructions[553] = {5'd1, 4'd2, 4'd4, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 33 {'a': 4, 'literal': 1, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 33, 'op': 'addl'}
    instructions[554] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 33 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 33, 'op': 'store'}
    instructions[555] = {5'd2, 4'd0, 4'd3, 16'd6};///tmp/tmpn6Oyv3/inline_c_file.c : 34 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 34, 'op': 'store'}
    instructions[556] = {5'd1, 4'd3, 4'd3, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 34 {'a': 3, 'literal': 1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 34, 'op': 'addl'}
    instructions[557] = {5'd2, 4'd0, 4'd3, 16'd7};///tmp/tmpn6Oyv3/inline_c_file.c : 34 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 34, 'op': 'store'}
    instructions[558] = {5'd1, 4'd3, 4'd3, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 34 {'a': 3, 'literal': 1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 34, 'op': 'addl'}
    instructions[559] = {5'd1, 4'd8, 4'd4, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 34 {'a': 4, 'literal': 1, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 34, 'op': 'addl'}
    instructions[560] = {5'd1, 4'd2, 4'd8, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 34 {'a': 8, 'literal': 0, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 34, 'op': 'addl'}
    instructions[561] = {5'd5, 4'd8, 4'd2, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 34 {'a': 2, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 34, 'op': 'load'}
    instructions[562] = {5'd2, 4'd0, 4'd3, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 34 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 34, 'op': 'store'}
    instructions[563] = {5'd1, 4'd3, 4'd3, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 34 {'a': 3, 'literal': 1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 34, 'op': 'addl'}
    instructions[564] = {5'd1, 4'd7, 4'd4, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 34 {'a': 4, 'literal': 0, 'z': 7, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 34, 'op': 'addl'}
    instructions[565] = {5'd1, 4'd4, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 34 {'a': 3, 'literal': 0, 'z': 4, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 34, 'op': 'addl'}
    instructions[566] = {5'd3, 4'd6, 4'd0, 16'd1079};///tmp/tmpn6Oyv3/inline_c_file.c : 34 {'z': 6, 'label': 1079, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 34, 'op': 'call'}
    instructions[567] = {5'd1, 4'd3, 4'd3, -16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 34 {'a': 3, 'literal': -1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 34, 'op': 'addl'}
    instructions[568] = {5'd1, 4'd3, 4'd3, -16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 34 {'a': 3, 'comment': 'pop', 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 34, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[569] = {5'd5, 4'd7, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 34 {'a': 3, 'z': 7, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 34, 'op': 'load'}
    instructions[570] = {5'd1, 4'd3, 4'd3, -16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 34 {'a': 3, 'comment': 'pop', 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 34, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[571] = {5'd5, 4'd6, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 34 {'a': 3, 'z': 6, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 34, 'op': 'load'}
    instructions[572] = {5'd1, 4'd3, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 34 {'a': 3, 'literal': 0, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 34, 'op': 'addl'}
    instructions[573] = {5'd2, 4'd0, 4'd3, 16'd6};///tmp/tmpn6Oyv3/inline_c_file.c : 34 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 34, 'op': 'store'}
    instructions[574] = {5'd1, 4'd3, 4'd3, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 34 {'a': 3, 'literal': 1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 34, 'op': 'addl'}
    instructions[575] = {5'd2, 4'd0, 4'd3, 16'd7};///tmp/tmpn6Oyv3/inline_c_file.c : 34 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 34, 'op': 'store'}
    instructions[576] = {5'd1, 4'd3, 4'd3, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 34 {'a': 3, 'literal': 1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 34, 'op': 'addl'}
    instructions[577] = {5'd0, 4'd8, 4'd0, 16'd31};///tmp/tmpn6Oyv3/inline_c_file.c : 35 {'literal': 31, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 35, 'op': 'literal'}
    instructions[578] = {5'd2, 4'd0, 4'd3, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 34 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 34, 'op': 'store'}
    instructions[579] = {5'd1, 4'd3, 4'd3, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 34 {'a': 3, 'literal': 1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 34, 'op': 'addl'}
    instructions[580] = {5'd1, 4'd7, 4'd4, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 34 {'a': 4, 'literal': 0, 'z': 7, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 34, 'op': 'addl'}
    instructions[581] = {5'd1, 4'd4, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 34 {'a': 3, 'literal': 0, 'z': 4, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 34, 'op': 'addl'}
    instructions[582] = {5'd3, 4'd6, 4'd0, 16'd687};///tmp/tmpn6Oyv3/inline_c_file.c : 34 {'z': 6, 'label': 687, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 34, 'op': 'call'}
    instructions[583] = {5'd1, 4'd3, 4'd3, -16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 34 {'a': 3, 'literal': -1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 34, 'op': 'addl'}
    instructions[584] = {5'd1, 4'd3, 4'd3, -16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 34 {'a': 3, 'comment': 'pop', 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 34, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[585] = {5'd5, 4'd7, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 34 {'a': 3, 'z': 7, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 34, 'op': 'load'}
    instructions[586] = {5'd1, 4'd3, 4'd3, -16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 34 {'a': 3, 'comment': 'pop', 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 34, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[587] = {5'd5, 4'd6, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 34 {'a': 3, 'z': 6, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 34, 'op': 'load'}
    instructions[588] = {5'd1, 4'd3, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 34 {'a': 3, 'literal': 0, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 34, 'op': 'addl'}
    instructions[589] = {5'd2, 4'd0, 4'd3, 16'd6};///tmp/tmpn6Oyv3/inline_c_file.c : 36 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 36, 'op': 'store'}
    instructions[590] = {5'd1, 4'd3, 4'd3, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 36 {'a': 3, 'literal': 1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 36, 'op': 'addl'}
    instructions[591] = {5'd2, 4'd0, 4'd3, 16'd7};///tmp/tmpn6Oyv3/inline_c_file.c : 36 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 36, 'op': 'store'}
    instructions[592] = {5'd1, 4'd3, 4'd3, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 36 {'a': 3, 'literal': 1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 36, 'op': 'addl'}
    instructions[593] = {5'd0, 4'd8, 4'd0, 16'd41};///tmp/tmpn6Oyv3/inline_c_file.c : 37 {'literal': 41, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 37, 'op': 'literal'}
    instructions[594] = {5'd2, 4'd0, 4'd3, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 36 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 36, 'op': 'store'}
    instructions[595] = {5'd1, 4'd3, 4'd3, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 36 {'a': 3, 'literal': 1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 36, 'op': 'addl'}
    instructions[596] = {5'd1, 4'd7, 4'd4, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 36 {'a': 4, 'literal': 0, 'z': 7, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 36, 'op': 'addl'}
    instructions[597] = {5'd1, 4'd4, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 36 {'a': 3, 'literal': 0, 'z': 4, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 36, 'op': 'addl'}
    instructions[598] = {5'd3, 4'd6, 4'd0, 16'd687};///tmp/tmpn6Oyv3/inline_c_file.c : 36 {'z': 6, 'label': 687, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 36, 'op': 'call'}
    instructions[599] = {5'd1, 4'd3, 4'd3, -16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 36 {'a': 3, 'literal': -1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 36, 'op': 'addl'}
    instructions[600] = {5'd1, 4'd3, 4'd3, -16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 36 {'a': 3, 'comment': 'pop', 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 36, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[601] = {5'd5, 4'd7, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 36 {'a': 3, 'z': 7, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 36, 'op': 'load'}
    instructions[602] = {5'd1, 4'd3, 4'd3, -16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 36 {'a': 3, 'comment': 'pop', 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 36, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[603] = {5'd5, 4'd6, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 36 {'a': 3, 'z': 6, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 36, 'op': 'load'}
    instructions[604] = {5'd1, 4'd3, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 36 {'a': 3, 'literal': 0, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 36, 'op': 'addl'}
    instructions[605] = {5'd2, 4'd0, 4'd3, 16'd6};///tmp/tmpn6Oyv3/inline_c_file.c : 38 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 38, 'op': 'store'}
    instructions[606] = {5'd1, 4'd3, 4'd3, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 38 {'a': 3, 'literal': 1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 38, 'op': 'addl'}
    instructions[607] = {5'd2, 4'd0, 4'd3, 16'd7};///tmp/tmpn6Oyv3/inline_c_file.c : 38 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 38, 'op': 'store'}
    instructions[608] = {5'd1, 4'd3, 4'd3, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 38 {'a': 3, 'literal': 1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 38, 'op': 'addl'}
    instructions[609] = {5'd1, 4'd7, 4'd4, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 38 {'a': 4, 'literal': 0, 'z': 7, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 38, 'op': 'addl'}
    instructions[610] = {5'd1, 4'd4, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 38 {'a': 3, 'literal': 0, 'z': 4, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 38, 'op': 'addl'}
    instructions[611] = {5'd3, 4'd6, 4'd0, 16'd778};///tmp/tmpn6Oyv3/inline_c_file.c : 38 {'z': 6, 'label': 778, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 38, 'op': 'call'}
    instructions[612] = {5'd1, 4'd3, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 38 {'a': 3, 'literal': 0, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 38, 'op': 'addl'}
    instructions[613] = {5'd1, 4'd3, 4'd3, -16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 38 {'a': 3, 'comment': 'pop', 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 38, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[614] = {5'd5, 4'd7, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 38 {'a': 3, 'z': 7, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 38, 'op': 'load'}
    instructions[615] = {5'd1, 4'd3, 4'd3, -16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 38 {'a': 3, 'comment': 'pop', 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 38, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[616] = {5'd5, 4'd6, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 38 {'a': 3, 'z': 6, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 38, 'op': 'load'}
    instructions[617] = {5'd0, 4'd2, 4'd0, 16'd37};///tmp/tmpn6Oyv3/inline_c_file.c : 38 {'literal': 37, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 38, 'op': 'literal'}
    instructions[618] = {5'd5, 4'd8, 4'd2, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 38 {'a': 2, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 38, 'op': 'load'}
    instructions[619] = {5'd1, 4'd2, 4'd4, 16'd2};///tmp/tmpn6Oyv3/inline_c_file.c : 38 {'a': 4, 'literal': 2, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 38, 'op': 'addl'}
    instructions[620] = {5'd2, 4'd0, 4'd2, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 38 {'a': 2, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 38, 'op': 'store'}
    instructions[621] = {5'd2, 4'd0, 4'd3, 16'd6};///tmp/tmpn6Oyv3/inline_c_file.c : 39 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 39, 'op': 'store'}
    instructions[622] = {5'd1, 4'd3, 4'd3, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 39 {'a': 3, 'literal': 1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 39, 'op': 'addl'}
    instructions[623] = {5'd2, 4'd0, 4'd3, 16'd7};///tmp/tmpn6Oyv3/inline_c_file.c : 39 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 39, 'op': 'store'}
    instructions[624] = {5'd1, 4'd3, 4'd3, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 39 {'a': 3, 'literal': 1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 39, 'op': 'addl'}
    instructions[625] = {5'd1, 4'd8, 4'd4, 16'd2};///tmp/tmpn6Oyv3/inline_c_file.c : 39 {'a': 4, 'literal': 2, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 39, 'op': 'addl'}
    instructions[626] = {5'd1, 4'd2, 4'd8, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 39 {'a': 8, 'literal': 0, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 39, 'op': 'addl'}
    instructions[627] = {5'd5, 4'd8, 4'd2, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 39 {'a': 2, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 39, 'op': 'load'}
    instructions[628] = {5'd2, 4'd0, 4'd3, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 39 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 39, 'op': 'store'}
    instructions[629] = {5'd1, 4'd3, 4'd3, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 39 {'a': 3, 'literal': 1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 39, 'op': 'addl'}
    instructions[630] = {5'd1, 4'd7, 4'd4, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 39 {'a': 4, 'literal': 0, 'z': 7, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 39, 'op': 'addl'}
    instructions[631] = {5'd1, 4'd4, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 39 {'a': 3, 'literal': 0, 'z': 4, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 39, 'op': 'addl'}
    instructions[632] = {5'd3, 4'd6, 4'd0, 16'd1079};///tmp/tmpn6Oyv3/inline_c_file.c : 39 {'z': 6, 'label': 1079, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 39, 'op': 'call'}
    instructions[633] = {5'd1, 4'd3, 4'd3, -16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 39 {'a': 3, 'literal': -1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 39, 'op': 'addl'}
    instructions[634] = {5'd1, 4'd3, 4'd3, -16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 39 {'a': 3, 'comment': 'pop', 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 39, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[635] = {5'd5, 4'd7, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 39 {'a': 3, 'z': 7, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 39, 'op': 'load'}
    instructions[636] = {5'd1, 4'd3, 4'd3, -16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 39 {'a': 3, 'comment': 'pop', 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 39, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[637] = {5'd5, 4'd6, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 39 {'a': 3, 'z': 6, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 39, 'op': 'load'}
    instructions[638] = {5'd1, 4'd3, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 39 {'a': 3, 'literal': 0, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 39, 'op': 'addl'}
    instructions[639] = {5'd2, 4'd0, 4'd3, 16'd6};///tmp/tmpn6Oyv3/inline_c_file.c : 39 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 39, 'op': 'store'}
    instructions[640] = {5'd1, 4'd3, 4'd3, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 39 {'a': 3, 'literal': 1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 39, 'op': 'addl'}
    instructions[641] = {5'd2, 4'd0, 4'd3, 16'd7};///tmp/tmpn6Oyv3/inline_c_file.c : 39 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 39, 'op': 'store'}
    instructions[642] = {5'd1, 4'd3, 4'd3, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 39 {'a': 3, 'literal': 1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 39, 'op': 'addl'}
    instructions[643] = {5'd0, 4'd8, 4'd0, 16'd108};///tmp/tmpn6Oyv3/inline_c_file.c : 40 {'literal': 108, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 40, 'op': 'literal'}
    instructions[644] = {5'd2, 4'd0, 4'd3, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 39 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 39, 'op': 'store'}
    instructions[645] = {5'd1, 4'd3, 4'd3, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 39 {'a': 3, 'literal': 1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 39, 'op': 'addl'}
    instructions[646] = {5'd1, 4'd7, 4'd4, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 39 {'a': 4, 'literal': 0, 'z': 7, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 39, 'op': 'addl'}
    instructions[647] = {5'd1, 4'd4, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 39 {'a': 3, 'literal': 0, 'z': 4, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 39, 'op': 'addl'}
    instructions[648] = {5'd3, 4'd6, 4'd0, 16'd687};///tmp/tmpn6Oyv3/inline_c_file.c : 39 {'z': 6, 'label': 687, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 39, 'op': 'call'}
    instructions[649] = {5'd1, 4'd3, 4'd3, -16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 39 {'a': 3, 'literal': -1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 39, 'op': 'addl'}
    instructions[650] = {5'd1, 4'd3, 4'd3, -16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 39 {'a': 3, 'comment': 'pop', 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 39, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[651] = {5'd5, 4'd7, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 39 {'a': 3, 'z': 7, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 39, 'op': 'load'}
    instructions[652] = {5'd1, 4'd3, 4'd3, -16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 39 {'a': 3, 'comment': 'pop', 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 39, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[653] = {5'd5, 4'd6, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 39 {'a': 3, 'z': 6, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 39, 'op': 'load'}
    instructions[654] = {5'd1, 4'd3, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 39 {'a': 3, 'literal': 0, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 39, 'op': 'addl'}
    instructions[655] = {5'd2, 4'd0, 4'd3, 16'd6};///tmp/tmpn6Oyv3/inline_c_file.c : 41 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 41, 'op': 'store'}
    instructions[656] = {5'd1, 4'd3, 4'd3, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 41 {'a': 3, 'literal': 1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 41, 'op': 'addl'}
    instructions[657] = {5'd2, 4'd0, 4'd3, 16'd7};///tmp/tmpn6Oyv3/inline_c_file.c : 41 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 41, 'op': 'store'}
    instructions[658] = {5'd1, 4'd3, 4'd3, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 41 {'a': 3, 'literal': 1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 41, 'op': 'addl'}
    instructions[659] = {5'd1, 4'd8, 4'd4, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 41 {'a': 4, 'literal': 0, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 41, 'op': 'addl'}
    instructions[660] = {5'd1, 4'd2, 4'd8, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 41 {'a': 8, 'literal': 0, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 41, 'op': 'addl'}
    instructions[661] = {5'd5, 4'd8, 4'd2, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 41 {'a': 2, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 41, 'op': 'load'}
    instructions[662] = {5'd2, 4'd0, 4'd3, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 41 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 41, 'op': 'store'}
    instructions[663] = {5'd1, 4'd3, 4'd3, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 41 {'a': 3, 'literal': 1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 41, 'op': 'addl'}
    instructions[664] = {5'd1, 4'd8, 4'd4, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 41 {'a': 4, 'literal': 1, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 41, 'op': 'addl'}
    instructions[665] = {5'd1, 4'd2, 4'd8, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 41 {'a': 8, 'literal': 0, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 41, 'op': 'addl'}
    instructions[666] = {5'd5, 4'd8, 4'd2, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 41 {'a': 2, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 41, 'op': 'load'}
    instructions[667] = {5'd2, 4'd0, 4'd3, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 41 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 41, 'op': 'store'}
    instructions[668] = {5'd1, 4'd3, 4'd3, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 41 {'a': 3, 'literal': 1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 41, 'op': 'addl'}
    instructions[669] = {5'd1, 4'd8, 4'd4, 16'd2};///tmp/tmpn6Oyv3/inline_c_file.c : 41 {'a': 4, 'literal': 2, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 41, 'op': 'addl'}
    instructions[670] = {5'd1, 4'd2, 4'd8, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 41 {'a': 8, 'literal': 0, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 41, 'op': 'addl'}
    instructions[671] = {5'd5, 4'd8, 4'd2, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 41 {'a': 2, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 41, 'op': 'load'}
    instructions[672] = {5'd2, 4'd0, 4'd3, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 41 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 41, 'op': 'store'}
    instructions[673] = {5'd1, 4'd3, 4'd3, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 41 {'a': 3, 'literal': 1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 41, 'op': 'addl'}
    instructions[674] = {5'd1, 4'd7, 4'd4, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 41 {'a': 4, 'literal': 0, 'z': 7, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 41, 'op': 'addl'}
    instructions[675] = {5'd1, 4'd4, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 41 {'a': 3, 'literal': 0, 'z': 4, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 41, 'op': 'addl'}
    instructions[676] = {5'd3, 4'd6, 4'd0, 16'd1235};///tmp/tmpn6Oyv3/inline_c_file.c : 41 {'z': 6, 'label': 1235, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 41, 'op': 'call'}
    instructions[677] = {5'd1, 4'd3, 4'd3, -16'd3};///tmp/tmpn6Oyv3/inline_c_file.c : 41 {'a': 3, 'literal': -3, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 41, 'op': 'addl'}
    instructions[678] = {5'd1, 4'd3, 4'd3, -16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 41 {'a': 3, 'comment': 'pop', 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 41, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[679] = {5'd5, 4'd7, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 41 {'a': 3, 'z': 7, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 41, 'op': 'load'}
    instructions[680] = {5'd1, 4'd3, 4'd3, -16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 41 {'a': 3, 'comment': 'pop', 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 41, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[681] = {5'd5, 4'd6, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 41 {'a': 3, 'z': 6, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 41, 'op': 'load'}
    instructions[682] = {5'd1, 4'd3, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 41 {'a': 3, 'literal': 0, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 41, 'op': 'addl'}
    instructions[683] = {5'd6, 4'd0, 4'd0, 16'd457};///tmp/tmpn6Oyv3/inline_c_file.c : 25 {'label': 457, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 25, 'op': 'goto'}
    instructions[684] = {5'd1, 4'd3, 4'd4, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 17 {'a': 4, 'literal': 0, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 17, 'op': 'addl'}
    instructions[685] = {5'd1, 4'd4, 4'd7, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 17 {'a': 7, 'literal': 0, 'z': 4, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 17, 'op': 'addl'}
    instructions[686] = {5'd7, 4'd0, 4'd6, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 17 {'a': 6, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 17, 'op': 'return'}
    instructions[687] = {5'd1, 4'd3, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73 {'a': 3, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73, 'op': 'addl'}
    instructions[688] = {5'd2, 4'd0, 4'd3, 16'd6};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'store'}
    instructions[689] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[690] = {5'd2, 4'd0, 4'd3, 16'd7};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'store'}
    instructions[691] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[692] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[693] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[694] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'load'}
    instructions[695] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'store'}
    instructions[696] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[697] = {5'd0, 4'd8, 4'd0, 16'd113};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'literal': 113, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'literal'}
    instructions[698] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[699] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'load'}
    instructions[700] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'store'}
    instructions[701] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[702] = {5'd1, 4'd7, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 4, 'literal': 0, 'z': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[703] = {5'd1, 4'd4, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[704] = {5'd3, 4'd6, 4'd0, 16'd714};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'z': 6, 'label': 714, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'call'}
    instructions[705] = {5'd1, 4'd3, 4'd3, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': -2, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[706] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[707] = {5'd5, 4'd7, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'z': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'load'}
    instructions[708] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[709] = {5'd5, 4'd6, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'z': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'load'}
    instructions[710] = {5'd1, 4'd3, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[711] = {5'd1, 4'd3, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73 {'a': 4, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73, 'op': 'addl'}
    instructions[712] = {5'd1, 4'd4, 4'd7, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73 {'a': 7, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73, 'op': 'addl'}
    instructions[713] = {5'd7, 4'd0, 4'd6, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73 {'a': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73, 'op': 'return'}
    instructions[714] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23, 'op': 'addl'}
    instructions[715] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 24 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 24, 'op': 'literal'}
    instructions[716] = {5'd1, 4'd2, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 24 {'a': 4, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 24, 'op': 'addl'}
    instructions[717] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 24 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 24, 'op': 'store'}
    instructions[718] = {5'd1, 4'd8, 4'd4, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 4, 'literal': -2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'addl'}
    instructions[719] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'addl'}
    instructions[720] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'load'}
    instructions[721] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'store'}
    instructions[722] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'addl'}
    instructions[723] = {5'd1, 4'd8, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 4, 'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'addl'}
    instructions[724] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'addl'}
    instructions[725] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'load'}
    instructions[726] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[727] = {5'd5, 4'd2, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 3, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'load'}
    instructions[728] = {5'd8, 4'd8, 4'd8, 16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 8, 'z': 8, 'b': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'add'}
    instructions[729] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'addl'}
    instructions[730] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'load'}
    instructions[731] = {5'd9, 4'd0, 4'd8, 16'd773};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 29 {'a': 8, 'label': 773, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 29, 'op': 'jmp_if_false'}
    instructions[732] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[733] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[734] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'load'}
    instructions[735] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'store'}
    instructions[736] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[737] = {5'd1, 4'd8, 4'd4, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 4, 'literal': -2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[738] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[739] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'load'}
    instructions[740] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'store'}
    instructions[741] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[742] = {5'd1, 4'd8, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 4, 'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[743] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[744] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'load'}
    instructions[745] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[746] = {5'd5, 4'd2, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'load'}
    instructions[747] = {5'd8, 4'd8, 4'd8, 16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 8, 'z': 8, 'b': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'add'}
    instructions[748] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[749] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'load'}
    instructions[750] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[751] = {5'd5, 4'd0, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'z': 0, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'load'}
    instructions[752] = {5'd10, 4'd0, 4'd0, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 0, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'write'}
    instructions[753] = {5'd1, 4'd3, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[754] = {5'd1, 4'd8, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 4, 'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[755] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[756] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'load'}
    instructions[757] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'store'}
    instructions[758] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[759] = {5'd0, 4'd8, 4'd0, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'literal': 1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'literal'}
    instructions[760] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'store'}
    instructions[761] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[762] = {5'd1, 4'd8, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 4, 'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[763] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[764] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'load'}
    instructions[765] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[766] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'load'}
    instructions[767] = {5'd8, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'add'}
    instructions[768] = {5'd1, 4'd2, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 4, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[769] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'store'}
    instructions[770] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[771] = {5'd5, 4'd8, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'load'}
    instructions[772] = {5'd6, 4'd0, 4'd0, 16'd774};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 29 {'label': 774, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 29, 'op': 'goto'}
    instructions[773] = {5'd6, 4'd0, 4'd0, 16'd775};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 29 {'label': 775, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 29, 'op': 'goto'}
    instructions[774] = {5'd6, 4'd0, 4'd0, 16'd718};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'label': 718, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'goto'}
    instructions[775] = {5'd1, 4'd3, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23 {'a': 4, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23, 'op': 'addl'}
    instructions[776] = {5'd1, 4'd4, 4'd7, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23 {'a': 7, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23, 'op': 'addl'}
    instructions[777] = {5'd7, 4'd0, 4'd6, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23 {'a': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23, 'op': 'return'}
    instructions[778] = {5'd1, 4'd3, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 151 {'a': 3, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 151, 'op': 'addl'}
    instructions[779] = {5'd2, 4'd0, 4'd3, 16'd6};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152, 'op': 'store'}
    instructions[780] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152, 'op': 'addl'}
    instructions[781] = {5'd2, 4'd0, 4'd3, 16'd7};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152, 'op': 'store'}
    instructions[782] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152, 'op': 'addl'}
    instructions[783] = {5'd0, 4'd8, 4'd0, 16'd38};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152 {'literal': 38, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152, 'op': 'literal'}
    instructions[784] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152, 'op': 'addl'}
    instructions[785] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152, 'op': 'load'}
    instructions[786] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152, 'op': 'store'}
    instructions[787] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152, 'op': 'addl'}
    instructions[788] = {5'd1, 4'd7, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152 {'a': 4, 'literal': 0, 'z': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152, 'op': 'addl'}
    instructions[789] = {5'd1, 4'd4, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152 {'a': 3, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152, 'op': 'addl'}
    instructions[790] = {5'd3, 4'd6, 4'd0, 16'd803};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152 {'z': 6, 'label': 803, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152, 'op': 'call'}
    instructions[791] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152 {'a': 3, 'literal': -1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152, 'op': 'addl'}
    instructions[792] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[793] = {5'd5, 4'd7, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152 {'a': 3, 'z': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152, 'op': 'load'}
    instructions[794] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[795] = {5'd5, 4'd6, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152 {'a': 3, 'z': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152, 'op': 'load'}
    instructions[796] = {5'd0, 4'd2, 4'd0, 16'd40};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152 {'literal': 40, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152, 'op': 'literal'}
    instructions[797] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152, 'op': 'load'}
    instructions[798] = {5'd0, 4'd2, 4'd0, 16'd37};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152 {'literal': 37, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152, 'op': 'literal'}
    instructions[799] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152, 'op': 'store'}
    instructions[800] = {5'd1, 4'd3, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152 {'a': 4, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152, 'op': 'addl'}
    instructions[801] = {5'd1, 4'd4, 4'd7, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152 {'a': 7, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152, 'op': 'addl'}
    instructions[802] = {5'd7, 4'd0, 4'd6, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152 {'a': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 152, 'op': 'return'}
    instructions[803] = {5'd1, 4'd3, 4'd3, 16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 13 {'a': 3, 'literal': 2, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 13, 'op': 'addl'}
    instructions[804] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 16 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 16, 'op': 'literal'}
    instructions[805] = {5'd1, 4'd2, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 16 {'a': 4, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 16, 'op': 'addl'}
    instructions[806] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 16 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 16, 'op': 'store'}
    instructions[807] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 18 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 18, 'op': 'addl'}
    instructions[808] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 18 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 18, 'op': 'addl'}
    instructions[809] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 18 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 18, 'op': 'load'}
    instructions[810] = {5'd11, 4'd8, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 18 {'a': 8, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 18, 'op': 'read'}
    instructions[811] = {5'd1, 4'd2, 4'd4, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 18 {'a': 4, 'literal': 1, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 18, 'op': 'addl'}
    instructions[812] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 18 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 18, 'op': 'store'}
    instructions[813] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19, 'op': 'literal'}
    instructions[814] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19, 'op': 'store'}
    instructions[815] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19, 'op': 'addl'}
    instructions[816] = {5'd2, 4'd0, 4'd3, 16'd6};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19, 'op': 'store'}
    instructions[817] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19, 'op': 'addl'}
    instructions[818] = {5'd2, 4'd0, 4'd3, 16'd7};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19, 'op': 'store'}
    instructions[819] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19, 'op': 'addl'}
    instructions[820] = {5'd1, 4'd8, 4'd4, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19 {'a': 4, 'literal': 1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19, 'op': 'addl'}
    instructions[821] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19, 'op': 'addl'}
    instructions[822] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19, 'op': 'load'}
    instructions[823] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19, 'op': 'store'}
    instructions[824] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19, 'op': 'addl'}
    instructions[825] = {5'd1, 4'd7, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19 {'a': 4, 'literal': 0, 'z': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19, 'op': 'addl'}
    instructions[826] = {5'd1, 4'd4, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19 {'a': 3, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19, 'op': 'addl'}
    instructions[827] = {5'd3, 4'd6, 4'd0, 16'd890};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19 {'z': 6, 'label': 890, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19, 'op': 'call'}
    instructions[828] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19 {'a': 3, 'literal': -1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19, 'op': 'addl'}
    instructions[829] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[830] = {5'd5, 4'd7, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19 {'a': 3, 'z': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19, 'op': 'load'}
    instructions[831] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[832] = {5'd5, 4'd6, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19 {'a': 3, 'z': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19, 'op': 'load'}
    instructions[833] = {5'd0, 4'd2, 4'd0, 16'd30};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19 {'literal': 30, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19, 'op': 'literal'}
    instructions[834] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19, 'op': 'load'}
    instructions[835] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[836] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19, 'op': 'load'}
    instructions[837] = {5'd12, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19, 'op': 'equal'}
    instructions[838] = {5'd9, 4'd0, 4'd8, 16'd841};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19 {'a': 8, 'label': 841, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19, 'op': 'jmp_if_false'}
    instructions[839] = {5'd6, 4'd0, 4'd0, 16'd882};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19 {'label': 882, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19, 'op': 'goto'}
    instructions[840] = {5'd6, 4'd0, 4'd0, 16'd841};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19 {'label': 841, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 19, 'op': 'goto'}
    instructions[841] = {5'd0, 4'd8, 4'd0, 16'd4};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 20 {'literal': 4, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 20, 'op': 'literal'}
    instructions[842] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 20 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 20, 'op': 'store'}
    instructions[843] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 20 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 20, 'op': 'addl'}
    instructions[844] = {5'd1, 4'd8, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 20 {'a': 4, 'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 20, 'op': 'addl'}
    instructions[845] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 20 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 20, 'op': 'addl'}
    instructions[846] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 20 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 20, 'op': 'load'}
    instructions[847] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 20 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 20, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[848] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 20 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 20, 'op': 'load'}
    instructions[849] = {5'd13, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 20 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 20, 'op': 'shift_left'}
    instructions[850] = {5'd1, 4'd2, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 20 {'a': 4, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 20, 'op': 'addl'}
    instructions[851] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 20 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 20, 'op': 'store'}
    instructions[852] = {5'd2, 4'd0, 4'd3, 16'd6};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21, 'op': 'store'}
    instructions[853] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21, 'op': 'addl'}
    instructions[854] = {5'd2, 4'd0, 4'd3, 16'd7};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21, 'op': 'store'}
    instructions[855] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21, 'op': 'addl'}
    instructions[856] = {5'd1, 4'd8, 4'd4, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21 {'a': 4, 'literal': 1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21, 'op': 'addl'}
    instructions[857] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21, 'op': 'addl'}
    instructions[858] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21, 'op': 'load'}
    instructions[859] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21, 'op': 'store'}
    instructions[860] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21, 'op': 'addl'}
    instructions[861] = {5'd1, 4'd7, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21 {'a': 4, 'literal': 0, 'z': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21, 'op': 'addl'}
    instructions[862] = {5'd1, 4'd4, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21 {'a': 3, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21, 'op': 'addl'}
    instructions[863] = {5'd3, 4'd6, 4'd0, 16'd955};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21 {'z': 6, 'label': 955, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21, 'op': 'call'}
    instructions[864] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21 {'a': 3, 'literal': -1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21, 'op': 'addl'}
    instructions[865] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[866] = {5'd5, 4'd7, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21 {'a': 3, 'z': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21, 'op': 'load'}
    instructions[867] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[868] = {5'd5, 4'd6, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21 {'a': 3, 'z': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21, 'op': 'load'}
    instructions[869] = {5'd0, 4'd2, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21 {'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21, 'op': 'literal'}
    instructions[870] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21, 'op': 'load'}
    instructions[871] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21, 'op': 'store'}
    instructions[872] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21, 'op': 'addl'}
    instructions[873] = {5'd1, 4'd8, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21 {'a': 4, 'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21, 'op': 'addl'}
    instructions[874] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21, 'op': 'addl'}
    instructions[875] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21, 'op': 'load'}
    instructions[876] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[877] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21, 'op': 'load'}
    instructions[878] = {5'd8, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21, 'op': 'add'}
    instructions[879] = {5'd1, 4'd2, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21 {'a': 4, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21, 'op': 'addl'}
    instructions[880] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 21, 'op': 'store'}
    instructions[881] = {5'd6, 4'd0, 4'd0, 16'd807};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 17 {'label': 807, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 17, 'op': 'goto'}
    instructions[882] = {5'd1, 4'd8, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 23 {'a': 4, 'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 23, 'op': 'addl'}
    instructions[883] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 23 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 23, 'op': 'addl'}
    instructions[884] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 23 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 23, 'op': 'load'}
    instructions[885] = {5'd0, 4'd2, 4'd0, 16'd40};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 23 {'literal': 40, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 23, 'op': 'literal'}
    instructions[886] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 23 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 23, 'op': 'store'}
    instructions[887] = {5'd1, 4'd3, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 23 {'a': 4, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 23, 'op': 'addl'}
    instructions[888] = {5'd1, 4'd4, 4'd7, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 23 {'a': 7, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 23, 'op': 'addl'}
    instructions[889] = {5'd7, 4'd0, 4'd6, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 23 {'a': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 23, 'op': 'return'}
    instructions[890] = {5'd1, 4'd3, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 240 {'a': 3, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 240, 'op': 'addl'}
    instructions[891] = {5'd0, 4'd8, 4'd0, 16'd65};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'literal': 65, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'literal'}
    instructions[892] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'store'}
    instructions[893] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'addl'}
    instructions[894] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'addl'}
    instructions[895] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'addl'}
    instructions[896] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'load'}
    instructions[897] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[898] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'load'}
    instructions[899] = {5'd14, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'greater_equal'}
    instructions[900] = {5'd9, 4'd0, 4'd8, 16'd910};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 8, 'label': 910, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'jmp_if_false'}
    instructions[901] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'addl'}
    instructions[902] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'addl'}
    instructions[903] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'load'}
    instructions[904] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'store'}
    instructions[905] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'addl'}
    instructions[906] = {5'd0, 4'd8, 4'd0, 16'd70};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'literal': 70, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'literal'}
    instructions[907] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[908] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'load'}
    instructions[909] = {5'd14, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'greater_equal'}
    instructions[910] = {5'd15, 4'd0, 4'd8, 16'd930};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 8, 'label': 930, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'jmp_if_true'}
    instructions[911] = {5'd0, 4'd8, 4'd0, 16'd97};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'literal': 97, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'literal'}
    instructions[912] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'store'}
    instructions[913] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'addl'}
    instructions[914] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'addl'}
    instructions[915] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'addl'}
    instructions[916] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'load'}
    instructions[917] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[918] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'load'}
    instructions[919] = {5'd14, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'greater_equal'}
    instructions[920] = {5'd9, 4'd0, 4'd8, 16'd930};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 8, 'label': 930, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'jmp_if_false'}
    instructions[921] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'addl'}
    instructions[922] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'addl'}
    instructions[923] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'load'}
    instructions[924] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'store'}
    instructions[925] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'addl'}
    instructions[926] = {5'd0, 4'd8, 4'd0, 16'd102};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'literal': 102, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'literal'}
    instructions[927] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[928] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'load'}
    instructions[929] = {5'd14, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'greater_equal'}
    instructions[930] = {5'd15, 4'd0, 4'd8, 16'd950};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 8, 'label': 950, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'jmp_if_true'}
    instructions[931] = {5'd0, 4'd8, 4'd0, 16'd48};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'literal': 48, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'literal'}
    instructions[932] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'store'}
    instructions[933] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'addl'}
    instructions[934] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'addl'}
    instructions[935] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'addl'}
    instructions[936] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'load'}
    instructions[937] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[938] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'load'}
    instructions[939] = {5'd14, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'greater_equal'}
    instructions[940] = {5'd9, 4'd0, 4'd8, 16'd950};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 8, 'label': 950, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'jmp_if_false'}
    instructions[941] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'addl'}
    instructions[942] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'addl'}
    instructions[943] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'load'}
    instructions[944] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'store'}
    instructions[945] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'addl'}
    instructions[946] = {5'd0, 4'd8, 4'd0, 16'd57};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'literal': 57, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'literal'}
    instructions[947] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[948] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'load'}
    instructions[949] = {5'd14, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'greater_equal'}
    instructions[950] = {5'd0, 4'd2, 4'd0, 16'd30};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'literal': 30, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'literal'}
    instructions[951] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'store'}
    instructions[952] = {5'd1, 4'd3, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 4, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'addl'}
    instructions[953] = {5'd1, 4'd4, 4'd7, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 7, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'addl'}
    instructions[954] = {5'd7, 4'd0, 4'd6, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241 {'a': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 241, 'op': 'return'}
    instructions[955] = {5'd1, 4'd3, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 6 {'a': 3, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 6, 'op': 'addl'}
    instructions[956] = {5'd0, 4'd8, 4'd0, 16'd48};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7 {'literal': 48, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7, 'op': 'literal'}
    instructions[957] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7, 'op': 'store'}
    instructions[958] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7, 'op': 'addl'}
    instructions[959] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7, 'op': 'addl'}
    instructions[960] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7, 'op': 'addl'}
    instructions[961] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7, 'op': 'load'}
    instructions[962] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[963] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7, 'op': 'load'}
    instructions[964] = {5'd14, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7, 'op': 'greater_equal'}
    instructions[965] = {5'd9, 4'd0, 4'd8, 16'd975};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7 {'a': 8, 'label': 975, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7, 'op': 'jmp_if_false'}
    instructions[966] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7, 'op': 'addl'}
    instructions[967] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7, 'op': 'addl'}
    instructions[968] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7, 'op': 'load'}
    instructions[969] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7, 'op': 'store'}
    instructions[970] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7, 'op': 'addl'}
    instructions[971] = {5'd0, 4'd8, 4'd0, 16'd57};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7 {'literal': 57, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7, 'op': 'literal'}
    instructions[972] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[973] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7, 'op': 'load'}
    instructions[974] = {5'd14, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7, 'op': 'greater_equal'}
    instructions[975] = {5'd9, 4'd0, 4'd8, 16'd991};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7 {'a': 8, 'label': 991, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7, 'op': 'jmp_if_false'}
    instructions[976] = {5'd0, 4'd8, 4'd0, 16'd48};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7 {'literal': 48, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7, 'op': 'literal'}
    instructions[977] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7, 'op': 'store'}
    instructions[978] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7, 'op': 'addl'}
    instructions[979] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7, 'op': 'addl'}
    instructions[980] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7, 'op': 'addl'}
    instructions[981] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7, 'op': 'load'}
    instructions[982] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[983] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7, 'op': 'load'}
    instructions[984] = {5'd16, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7, 'op': 'subtract'}
    instructions[985] = {5'd0, 4'd2, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7 {'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7, 'op': 'literal'}
    instructions[986] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7, 'op': 'store'}
    instructions[987] = {5'd1, 4'd3, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7 {'a': 4, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7, 'op': 'addl'}
    instructions[988] = {5'd1, 4'd4, 4'd7, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7 {'a': 7, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7, 'op': 'addl'}
    instructions[989] = {5'd7, 4'd0, 4'd6, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7 {'a': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7, 'op': 'return'}
    instructions[990] = {5'd6, 4'd0, 4'd0, 16'd991};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7 {'label': 991, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 7, 'op': 'goto'}
    instructions[991] = {5'd0, 4'd8, 4'd0, 16'd97};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8 {'literal': 97, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8, 'op': 'literal'}
    instructions[992] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8, 'op': 'store'}
    instructions[993] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8, 'op': 'addl'}
    instructions[994] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8, 'op': 'addl'}
    instructions[995] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8, 'op': 'addl'}
    instructions[996] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8, 'op': 'load'}
    instructions[997] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[998] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8, 'op': 'load'}
    instructions[999] = {5'd14, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8, 'op': 'greater_equal'}
    instructions[1000] = {5'd9, 4'd0, 4'd8, 16'd1010};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8 {'a': 8, 'label': 1010, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8, 'op': 'jmp_if_false'}
    instructions[1001] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8, 'op': 'addl'}
    instructions[1002] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8, 'op': 'addl'}
    instructions[1003] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8, 'op': 'load'}
    instructions[1004] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8, 'op': 'store'}
    instructions[1005] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8, 'op': 'addl'}
    instructions[1006] = {5'd0, 4'd8, 4'd0, 16'd102};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8 {'literal': 102, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8, 'op': 'literal'}
    instructions[1007] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1008] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8, 'op': 'load'}
    instructions[1009] = {5'd14, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8, 'op': 'greater_equal'}
    instructions[1010] = {5'd9, 4'd0, 4'd8, 16'd1032};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8 {'a': 8, 'label': 1032, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8, 'op': 'jmp_if_false'}
    instructions[1011] = {5'd0, 4'd8, 4'd0, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8 {'literal': 10, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8, 'op': 'literal'}
    instructions[1012] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8, 'op': 'store'}
    instructions[1013] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8, 'op': 'addl'}
    instructions[1014] = {5'd0, 4'd8, 4'd0, 16'd97};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8 {'literal': 97, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8, 'op': 'literal'}
    instructions[1015] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8, 'op': 'store'}
    instructions[1016] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8, 'op': 'addl'}
    instructions[1017] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8, 'op': 'addl'}
    instructions[1018] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8, 'op': 'addl'}
    instructions[1019] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8, 'op': 'load'}
    instructions[1020] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1021] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8, 'op': 'load'}
    instructions[1022] = {5'd16, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8, 'op': 'subtract'}
    instructions[1023] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1024] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8, 'op': 'load'}
    instructions[1025] = {5'd8, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8, 'op': 'add'}
    instructions[1026] = {5'd0, 4'd2, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8 {'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8, 'op': 'literal'}
    instructions[1027] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8, 'op': 'store'}
    instructions[1028] = {5'd1, 4'd3, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8 {'a': 4, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8, 'op': 'addl'}
    instructions[1029] = {5'd1, 4'd4, 4'd7, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8 {'a': 7, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8, 'op': 'addl'}
    instructions[1030] = {5'd7, 4'd0, 4'd6, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8 {'a': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8, 'op': 'return'}
    instructions[1031] = {5'd6, 4'd0, 4'd0, 16'd1032};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8 {'label': 1032, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 8, 'op': 'goto'}
    instructions[1032] = {5'd0, 4'd8, 4'd0, 16'd65};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9 {'literal': 65, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9, 'op': 'literal'}
    instructions[1033] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9, 'op': 'store'}
    instructions[1034] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9, 'op': 'addl'}
    instructions[1035] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9, 'op': 'addl'}
    instructions[1036] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9, 'op': 'addl'}
    instructions[1037] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9, 'op': 'load'}
    instructions[1038] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1039] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9, 'op': 'load'}
    instructions[1040] = {5'd14, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9, 'op': 'greater_equal'}
    instructions[1041] = {5'd9, 4'd0, 4'd8, 16'd1051};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9 {'a': 8, 'label': 1051, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9, 'op': 'jmp_if_false'}
    instructions[1042] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9, 'op': 'addl'}
    instructions[1043] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9, 'op': 'addl'}
    instructions[1044] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9, 'op': 'load'}
    instructions[1045] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9, 'op': 'store'}
    instructions[1046] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9, 'op': 'addl'}
    instructions[1047] = {5'd0, 4'd8, 4'd0, 16'd70};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9 {'literal': 70, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9, 'op': 'literal'}
    instructions[1048] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1049] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9, 'op': 'load'}
    instructions[1050] = {5'd14, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9, 'op': 'greater_equal'}
    instructions[1051] = {5'd9, 4'd0, 4'd8, 16'd1073};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9 {'a': 8, 'label': 1073, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9, 'op': 'jmp_if_false'}
    instructions[1052] = {5'd0, 4'd8, 4'd0, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9 {'literal': 10, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9, 'op': 'literal'}
    instructions[1053] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9, 'op': 'store'}
    instructions[1054] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9, 'op': 'addl'}
    instructions[1055] = {5'd0, 4'd8, 4'd0, 16'd65};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9 {'literal': 65, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9, 'op': 'literal'}
    instructions[1056] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9, 'op': 'store'}
    instructions[1057] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9, 'op': 'addl'}
    instructions[1058] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9, 'op': 'addl'}
    instructions[1059] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9, 'op': 'addl'}
    instructions[1060] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9, 'op': 'load'}
    instructions[1061] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1062] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9, 'op': 'load'}
    instructions[1063] = {5'd16, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9, 'op': 'subtract'}
    instructions[1064] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1065] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9, 'op': 'load'}
    instructions[1066] = {5'd8, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9, 'op': 'add'}
    instructions[1067] = {5'd0, 4'd2, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9 {'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9, 'op': 'literal'}
    instructions[1068] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9, 'op': 'store'}
    instructions[1069] = {5'd1, 4'd3, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9 {'a': 4, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9, 'op': 'addl'}
    instructions[1070] = {5'd1, 4'd4, 4'd7, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9 {'a': 7, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9, 'op': 'addl'}
    instructions[1071] = {5'd7, 4'd0, 4'd6, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9 {'a': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9, 'op': 'return'}
    instructions[1072] = {5'd6, 4'd0, 4'd0, 16'd1073};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9 {'label': 1073, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 9, 'op': 'goto'}
    instructions[1073] = {5'd0, 4'd8, 4'd0, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 10 {'literal': 10, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 10, 'op': 'literal'}
    instructions[1074] = {5'd0, 4'd2, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 10 {'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 10, 'op': 'literal'}
    instructions[1075] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 10 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 10, 'op': 'store'}
    instructions[1076] = {5'd1, 4'd3, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 10 {'a': 4, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 10, 'op': 'addl'}
    instructions[1077] = {5'd1, 4'd4, 4'd7, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 10 {'a': 7, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 10, 'op': 'addl'}
    instructions[1078] = {5'd7, 4'd0, 4'd6, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 10 {'a': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 10, 'op': 'return'}
    instructions[1079] = {5'd1, 4'd3, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 149 {'a': 3, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 149, 'op': 'addl'}
    instructions[1080] = {5'd2, 4'd0, 4'd3, 16'd6};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 150 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 150, 'op': 'store'}
    instructions[1081] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 150 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 150, 'op': 'addl'}
    instructions[1082] = {5'd2, 4'd0, 4'd3, 16'd7};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 150 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 150, 'op': 'store'}
    instructions[1083] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 150 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 150, 'op': 'addl'}
    instructions[1084] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 150 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 150, 'op': 'addl'}
    instructions[1085] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 150 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 150, 'op': 'addl'}
    instructions[1086] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 150 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 150, 'op': 'load'}
    instructions[1087] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 150 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 150, 'op': 'store'}
    instructions[1088] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 150 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 150, 'op': 'addl'}
    instructions[1089] = {5'd0, 4'd8, 4'd0, 16'd113};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 150 {'literal': 113, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 150, 'op': 'literal'}
    instructions[1090] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 150 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 150, 'op': 'addl'}
    instructions[1091] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 150 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 150, 'op': 'load'}
    instructions[1092] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 150 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 150, 'op': 'store'}
    instructions[1093] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 150 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 150, 'op': 'addl'}
    instructions[1094] = {5'd1, 4'd7, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 150 {'a': 4, 'literal': 0, 'z': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 150, 'op': 'addl'}
    instructions[1095] = {5'd1, 4'd4, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 150 {'a': 3, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 150, 'op': 'addl'}
    instructions[1096] = {5'd3, 4'd6, 4'd0, 16'd1106};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 150 {'z': 6, 'label': 1106, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 150, 'op': 'call'}
    instructions[1097] = {5'd1, 4'd3, 4'd3, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 150 {'a': 3, 'literal': -2, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 150, 'op': 'addl'}
    instructions[1098] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 150 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 150, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1099] = {5'd5, 4'd7, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 150 {'a': 3, 'z': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 150, 'op': 'load'}
    instructions[1100] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 150 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 150, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1101] = {5'd5, 4'd6, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 150 {'a': 3, 'z': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 150, 'op': 'load'}
    instructions[1102] = {5'd1, 4'd3, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 150 {'a': 3, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 150, 'op': 'addl'}
    instructions[1103] = {5'd1, 4'd3, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 149 {'a': 4, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 149, 'op': 'addl'}
    instructions[1104] = {5'd1, 4'd4, 4'd7, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 149 {'a': 7, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 149, 'op': 'addl'}
    instructions[1105] = {5'd7, 4'd0, 4'd6, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 149 {'a': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 149, 'op': 'return'}
    instructions[1106] = {5'd1, 4'd3, 4'd3, 16'd19};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 4 {'a': 3, 'literal': 19, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 4, 'op': 'addl'}
    instructions[1107] = {5'd0, 4'd8, 4'd0, 16'd48};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'literal': 48, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'literal'}
    instructions[1108] = {5'd1, 4'd2, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'a': 4, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'addl'}
    instructions[1109] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'store'}
    instructions[1110] = {5'd0, 4'd8, 4'd0, 16'd49};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'literal': 49, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'literal'}
    instructions[1111] = {5'd1, 4'd2, 4'd4, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'a': 4, 'literal': 1, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'addl'}
    instructions[1112] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'store'}
    instructions[1113] = {5'd0, 4'd8, 4'd0, 16'd50};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'literal': 50, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'literal'}
    instructions[1114] = {5'd1, 4'd2, 4'd4, 16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'a': 4, 'literal': 2, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'addl'}
    instructions[1115] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'store'}
    instructions[1116] = {5'd0, 4'd8, 4'd0, 16'd51};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'literal': 51, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'literal'}
    instructions[1117] = {5'd1, 4'd2, 4'd4, 16'd3};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'a': 4, 'literal': 3, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'addl'}
    instructions[1118] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'store'}
    instructions[1119] = {5'd0, 4'd8, 4'd0, 16'd52};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'literal': 52, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'literal'}
    instructions[1120] = {5'd1, 4'd2, 4'd4, 16'd4};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'a': 4, 'literal': 4, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'addl'}
    instructions[1121] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'store'}
    instructions[1122] = {5'd0, 4'd8, 4'd0, 16'd53};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'literal': 53, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'literal'}
    instructions[1123] = {5'd1, 4'd2, 4'd4, 16'd5};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'a': 4, 'literal': 5, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'addl'}
    instructions[1124] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'store'}
    instructions[1125] = {5'd0, 4'd8, 4'd0, 16'd54};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'literal': 54, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'literal'}
    instructions[1126] = {5'd1, 4'd2, 4'd4, 16'd6};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'a': 4, 'literal': 6, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'addl'}
    instructions[1127] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'store'}
    instructions[1128] = {5'd0, 4'd8, 4'd0, 16'd55};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'literal': 55, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'literal'}
    instructions[1129] = {5'd1, 4'd2, 4'd4, 16'd7};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'a': 4, 'literal': 7, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'addl'}
    instructions[1130] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'store'}
    instructions[1131] = {5'd0, 4'd8, 4'd0, 16'd56};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'literal': 56, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'literal'}
    instructions[1132] = {5'd1, 4'd2, 4'd4, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'a': 4, 'literal': 8, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'addl'}
    instructions[1133] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'store'}
    instructions[1134] = {5'd0, 4'd8, 4'd0, 16'd57};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'literal': 57, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'literal'}
    instructions[1135] = {5'd1, 4'd2, 4'd4, 16'd9};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'a': 4, 'literal': 9, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'addl'}
    instructions[1136] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'store'}
    instructions[1137] = {5'd0, 4'd8, 4'd0, 16'd97};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'literal': 97, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'literal'}
    instructions[1138] = {5'd1, 4'd2, 4'd4, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'a': 4, 'literal': 10, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'addl'}
    instructions[1139] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'store'}
    instructions[1140] = {5'd0, 4'd8, 4'd0, 16'd98};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'literal': 98, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'literal'}
    instructions[1141] = {5'd1, 4'd2, 4'd4, 16'd11};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'a': 4, 'literal': 11, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'addl'}
    instructions[1142] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'store'}
    instructions[1143] = {5'd0, 4'd8, 4'd0, 16'd99};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'literal': 99, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'literal'}
    instructions[1144] = {5'd1, 4'd2, 4'd4, 16'd12};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'a': 4, 'literal': 12, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'addl'}
    instructions[1145] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'store'}
    instructions[1146] = {5'd0, 4'd8, 4'd0, 16'd100};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'literal': 100, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'literal'}
    instructions[1147] = {5'd1, 4'd2, 4'd4, 16'd13};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'a': 4, 'literal': 13, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'addl'}
    instructions[1148] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'store'}
    instructions[1149] = {5'd0, 4'd8, 4'd0, 16'd101};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'literal': 101, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'literal'}
    instructions[1150] = {5'd1, 4'd2, 4'd4, 16'd14};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'a': 4, 'literal': 14, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'addl'}
    instructions[1151] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'store'}
    instructions[1152] = {5'd0, 4'd8, 4'd0, 16'd102};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'literal': 102, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'literal'}
    instructions[1153] = {5'd1, 4'd2, 4'd4, 16'd15};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'a': 4, 'literal': 15, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'addl'}
    instructions[1154] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'store'}
    instructions[1155] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'literal'}
    instructions[1156] = {5'd1, 4'd2, 4'd4, 16'd16};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'a': 4, 'literal': 16, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'addl'}
    instructions[1157] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 5, 'op': 'store'}
    instructions[1158] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7, 'op': 'literal'}
    instructions[1159] = {5'd1, 4'd2, 4'd4, 16'd17};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7 {'a': 4, 'literal': 17, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7, 'op': 'addl'}
    instructions[1160] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7, 'op': 'store'}
    instructions[1161] = {5'd1, 4'd8, 4'd4, 16'd17};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7 {'a': 4, 'literal': 17, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7, 'op': 'addl'}
    instructions[1162] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7, 'op': 'addl'}
    instructions[1163] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7, 'op': 'load'}
    instructions[1164] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7, 'op': 'store'}
    instructions[1165] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7, 'op': 'addl'}
    instructions[1166] = {5'd0, 4'd8, 4'd0, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7 {'literal': 8, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7, 'op': 'literal'}
    instructions[1167] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1168] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7, 'op': 'load'}
    instructions[1169] = {5'd17, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7, 'op': 'unsigned_greater'}
    instructions[1170] = {5'd9, 4'd0, 4'd8, 16'd1232};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7 {'a': 8, 'label': 1232, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7, 'op': 'jmp_if_false'}
    instructions[1171] = {5'd0, 4'd8, 4'd0, 16'd28};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 8 {'literal': 28, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 8, 'op': 'literal'}
    instructions[1172] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 8 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 8, 'op': 'store'}
    instructions[1173] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 8 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 8, 'op': 'addl'}
    instructions[1174] = {5'd1, 4'd8, 4'd4, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 8 {'a': 4, 'literal': -2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 8, 'op': 'addl'}
    instructions[1175] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 8 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 8, 'op': 'addl'}
    instructions[1176] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 8 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 8, 'op': 'load'}
    instructions[1177] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 8 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 8, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1178] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 8 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 8, 'op': 'load'}
    instructions[1179] = {5'd18, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 8 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 8, 'op': 'unsigned_shift_right'}
    instructions[1180] = {5'd1, 4'd2, 4'd4, 16'd18};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 8 {'a': 4, 'literal': 18, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 8, 'op': 'addl'}
    instructions[1181] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 8 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 8, 'op': 'store'}
    instructions[1182] = {5'd0, 4'd8, 4'd0, 16'd4};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 9 {'literal': 4, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 9, 'op': 'literal'}
    instructions[1183] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 9 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 9, 'op': 'store'}
    instructions[1184] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 9 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 9, 'op': 'addl'}
    instructions[1185] = {5'd1, 4'd8, 4'd4, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 9 {'a': 4, 'literal': -2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 9, 'op': 'addl'}
    instructions[1186] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 9 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 9, 'op': 'addl'}
    instructions[1187] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 9 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 9, 'op': 'load'}
    instructions[1188] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 9 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 9, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1189] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 9 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 9, 'op': 'load'}
    instructions[1190] = {5'd13, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 9 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 9, 'op': 'shift_left'}
    instructions[1191] = {5'd1, 4'd2, 4'd4, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 9 {'a': 4, 'literal': -2, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 9, 'op': 'addl'}
    instructions[1192] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 9 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 9, 'op': 'store'}
    instructions[1193] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 10 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 10, 'op': 'addl'}
    instructions[1194] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 10 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 10, 'op': 'addl'}
    instructions[1195] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 10 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 10, 'op': 'load'}
    instructions[1196] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 10 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 10, 'op': 'store'}
    instructions[1197] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 10 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 10, 'op': 'addl'}
    instructions[1198] = {5'd1, 4'd8, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 10 {'a': 4, 'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 10, 'op': 'addl'}
    instructions[1199] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 10 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 10, 'op': 'store'}
    instructions[1200] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 10 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 10, 'op': 'addl'}
    instructions[1201] = {5'd1, 4'd8, 4'd4, 16'd18};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 10 {'a': 4, 'literal': 18, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 10, 'op': 'addl'}
    instructions[1202] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 10 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 10, 'op': 'addl'}
    instructions[1203] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 10 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 10, 'op': 'load'}
    instructions[1204] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 10 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 10, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1205] = {5'd5, 4'd2, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 10 {'a': 3, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 10, 'op': 'load'}
    instructions[1206] = {5'd8, 4'd8, 4'd8, 16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 10 {'a': 8, 'z': 8, 'b': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 10, 'op': 'add'}
    instructions[1207] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 10 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 10, 'op': 'addl'}
    instructions[1208] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 10 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 10, 'op': 'load'}
    instructions[1209] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 10 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 10, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1210] = {5'd5, 4'd0, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 10 {'a': 3, 'z': 0, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 10, 'op': 'load'}
    instructions[1211] = {5'd10, 4'd0, 4'd0, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 10 {'a': 0, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 10, 'op': 'write'}
    instructions[1212] = {5'd1, 4'd3, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 10 {'a': 3, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 10, 'op': 'addl'}
    instructions[1213] = {5'd1, 4'd8, 4'd4, 16'd17};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7 {'a': 4, 'literal': 17, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7, 'op': 'addl'}
    instructions[1214] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7, 'op': 'addl'}
    instructions[1215] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7, 'op': 'load'}
    instructions[1216] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7, 'op': 'store'}
    instructions[1217] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7, 'op': 'addl'}
    instructions[1218] = {5'd0, 4'd8, 4'd0, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7 {'literal': 1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7, 'op': 'literal'}
    instructions[1219] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7, 'op': 'store'}
    instructions[1220] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7, 'op': 'addl'}
    instructions[1221] = {5'd1, 4'd8, 4'd4, 16'd17};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7 {'a': 4, 'literal': 17, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7, 'op': 'addl'}
    instructions[1222] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7, 'op': 'addl'}
    instructions[1223] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7, 'op': 'load'}
    instructions[1224] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1225] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7, 'op': 'load'}
    instructions[1226] = {5'd8, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7, 'op': 'add'}
    instructions[1227] = {5'd1, 4'd2, 4'd4, 16'd17};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7 {'a': 4, 'literal': 17, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7, 'op': 'addl'}
    instructions[1228] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7, 'op': 'store'}
    instructions[1229] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1230] = {5'd5, 4'd8, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7 {'a': 3, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7, 'op': 'load'}
    instructions[1231] = {5'd6, 4'd0, 4'd0, 16'd1161};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7 {'label': 1161, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 7, 'op': 'goto'}
    instructions[1232] = {5'd1, 4'd3, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 4 {'a': 4, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 4, 'op': 'addl'}
    instructions[1233] = {5'd1, 4'd4, 4'd7, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 4 {'a': 7, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 4, 'op': 'addl'}
    instructions[1234] = {5'd7, 4'd0, 4'd6, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 4 {'a': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 4, 'op': 'return'}
    instructions[1235] = {5'd1, 4'd3, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 11 {'a': 3, 'literal': 0, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 11, 'op': 'addl'}
    instructions[1236] = {5'd0, 4'd8, 4'd0, 16'd39};///tmp/tmpn6Oyv3/inline_c_file.c : 12 {'literal': 39, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 12, 'op': 'literal'}
    instructions[1237] = {5'd1, 4'd2, 4'd8, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 12 {'a': 8, 'literal': 0, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 12, 'op': 'addl'}
    instructions[1238] = {5'd5, 4'd8, 4'd2, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 12 {'a': 2, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 12, 'op': 'load'}
    instructions[1239] = {5'd2, 4'd0, 4'd3, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 12 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 12, 'op': 'store'}
    instructions[1240] = {5'd1, 4'd3, 4'd3, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 12 {'a': 3, 'literal': 1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 12, 'op': 'addl'}
    instructions[1241] = {5'd1, 4'd8, 4'd4, -16'd3};///tmp/tmpn6Oyv3/inline_c_file.c : 12 {'a': 4, 'literal': -3, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 12, 'op': 'addl'}
    instructions[1242] = {5'd1, 4'd2, 4'd8, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 12 {'a': 8, 'literal': 0, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 12, 'op': 'addl'}
    instructions[1243] = {5'd5, 4'd8, 4'd2, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 12 {'a': 2, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 12, 'op': 'load'}
    instructions[1244] = {5'd1, 4'd3, 4'd3, -16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 12 {'a': 3, 'comment': 'pop', 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 12, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1245] = {5'd5, 4'd0, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 12 {'a': 3, 'z': 0, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 12, 'op': 'load'}
    instructions[1246] = {5'd10, 4'd0, 4'd0, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 12 {'a': 0, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 12, 'op': 'write'}
    instructions[1247] = {5'd1, 4'd3, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 12 {'a': 3, 'literal': 0, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 12, 'op': 'addl'}
    instructions[1248] = {5'd0, 4'd8, 4'd0, 16'd106};///tmp/tmpn6Oyv3/inline_c_file.c : 13 {'literal': 106, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 13, 'op': 'literal'}
    instructions[1249] = {5'd1, 4'd2, 4'd8, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 13 {'a': 8, 'literal': 0, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 13, 'op': 'addl'}
    instructions[1250] = {5'd5, 4'd8, 4'd2, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 13 {'a': 2, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 13, 'op': 'load'}
    instructions[1251] = {5'd2, 4'd0, 4'd3, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 13 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 13, 'op': 'store'}
    instructions[1252] = {5'd1, 4'd3, 4'd3, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 13 {'a': 3, 'literal': 1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 13, 'op': 'addl'}
    instructions[1253] = {5'd1, 4'd8, 4'd4, -16'd2};///tmp/tmpn6Oyv3/inline_c_file.c : 13 {'a': 4, 'literal': -2, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 13, 'op': 'addl'}
    instructions[1254] = {5'd1, 4'd2, 4'd8, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 13 {'a': 8, 'literal': 0, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 13, 'op': 'addl'}
    instructions[1255] = {5'd5, 4'd8, 4'd2, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 13 {'a': 2, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 13, 'op': 'load'}
    instructions[1256] = {5'd1, 4'd3, 4'd3, -16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 13 {'a': 3, 'comment': 'pop', 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 13, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1257] = {5'd5, 4'd0, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 13 {'a': 3, 'z': 0, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 13, 'op': 'load'}
    instructions[1258] = {5'd10, 4'd0, 4'd0, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 13 {'a': 0, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 13, 'op': 'write'}
    instructions[1259] = {5'd1, 4'd3, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 13 {'a': 3, 'literal': 0, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 13, 'op': 'addl'}
    instructions[1260] = {5'd0, 4'd8, 4'd0, 16'd107};///tmp/tmpn6Oyv3/inline_c_file.c : 14 {'literal': 107, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 14, 'op': 'literal'}
    instructions[1261] = {5'd1, 4'd2, 4'd8, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 14 {'a': 8, 'literal': 0, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 14, 'op': 'addl'}
    instructions[1262] = {5'd5, 4'd8, 4'd2, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 14 {'a': 2, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 14, 'op': 'load'}
    instructions[1263] = {5'd2, 4'd0, 4'd3, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 14 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 14, 'op': 'store'}
    instructions[1264] = {5'd1, 4'd3, 4'd3, 16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 14 {'a': 3, 'literal': 1, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 14, 'op': 'addl'}
    instructions[1265] = {5'd1, 4'd8, 4'd4, -16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 14 {'a': 4, 'literal': -1, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 14, 'op': 'addl'}
    instructions[1266] = {5'd1, 4'd2, 4'd8, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 14 {'a': 8, 'literal': 0, 'z': 2, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 14, 'op': 'addl'}
    instructions[1267] = {5'd5, 4'd8, 4'd2, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 14 {'a': 2, 'z': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 14, 'op': 'load'}
    instructions[1268] = {5'd1, 4'd3, 4'd3, -16'd1};///tmp/tmpn6Oyv3/inline_c_file.c : 14 {'a': 3, 'comment': 'pop', 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 14, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1269] = {5'd5, 4'd0, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 14 {'a': 3, 'z': 0, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 14, 'op': 'load'}
    instructions[1270] = {5'd10, 4'd0, 4'd0, 16'd8};///tmp/tmpn6Oyv3/inline_c_file.c : 14 {'a': 0, 'b': 8, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 14, 'op': 'write'}
    instructions[1271] = {5'd1, 4'd3, 4'd3, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 14 {'a': 3, 'literal': 0, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 14, 'op': 'addl'}
    instructions[1272] = {5'd1, 4'd3, 4'd4, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 11 {'a': 4, 'literal': 0, 'z': 3, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 11, 'op': 'addl'}
    instructions[1273] = {5'd1, 4'd4, 4'd7, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 11 {'a': 7, 'literal': 0, 'z': 4, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 11, 'op': 'addl'}
    instructions[1274] = {5'd7, 4'd0, 4'd6, 16'd0};///tmp/tmpn6Oyv3/inline_c_file.c : 11 {'a': 6, 'trace': /tmp/tmpn6Oyv3/inline_c_file.c : 11, 'op': 'return'}
  end

  
  always @(posedge clk)
  begin
    load_data <= memory[load_address];
    if(store_enable && state == execute) begin
      memory[store_address] <= store_data;
    end
  end


  //////////////////////////////////////////////////////////////////////////////
  // PIPELINE STAGE 1 -- FETCH INSTRUCTION
  //                                                                            
  
  always @(posedge clk)
  begin
    //implement memory for instructions
    if (state == instruction_fetch || state == operand_fetch || state == execute) begin
      instruction <= instructions[program_counter];
      program_counter_1 <= program_counter;
    end
  end

  assign opcode    = instruction[28:24];
  assign address_z = instruction[23:20];
  assign address_a = instruction[19:16];
  assign address_b = instruction[3:0];
  assign literal   = instruction[15:0];

  //////////////////////////////////////////////////////////////////////////////
  // PIPELINE STAGE 2 -- FETCH OPERANDS
  //                                                                            
  
  always @(posedge clk)
  begin
    if (write_enable) begin
      registers[address_z_3] <= result;
    end
    if (state == operand_fetch || state == execute) begin
      opcode_2 <= opcode;
      literal_2 <= literal;
      address_a_2 <= address_a;
      address_b_2 <= address_b;
      address_z_2 <= address_z;
      program_counter_2 <= program_counter_1;
    end
  end
  assign register_a = registers[address_a_2];
  assign register_b = registers[address_b_2];
  assign operand_a = (address_a_2 == address_z_3 && write_enable)?result:register_a;
  assign operand_b = (address_b_2 == address_z_3 && write_enable)?result:register_b;
  assign store_address = operand_a;
  assign load_address = operand_a;
  assign store_data = operand_b;
  assign store_enable = (opcode_2==2);

  //////////////////////////////////////////////////////////////////////////////
  // PIPELINE STAGE 3 -- EXECUTE
  //                                                                            
  
  always @(posedge clk)
  begin

  write_enable <= 0;
  timer_clock <= timer_clock + 1;
  case(state)

    //instruction_fetch
    instruction_fetch: begin
      program_counter <= program_counter + 1;
      state <= operand_fetch;
    end
    //operand_fetch
    operand_fetch: begin
      program_counter <= program_counter + 1;
      state <= execute;
    end
    //execute
    execute: begin
      program_counter <= program_counter + 1;
      address_z_3 <= address_z_2;
      case(opcode_2)

        //literal
        16'd0:
        begin
          result<=$signed(literal_2);
          write_enable <= 1;
        end

        //addl
        16'd1:
        begin
          result<=operand_a + literal_2;
          write_enable <= 1;
        end

        //store
        16'd2:
        begin
        end

        //call
        16'd3:
        begin
          result <= program_counter_2 + 1;
          write_enable <= 1;
          program_counter <= literal_2;
          state <= instruction_fetch;
        end

        //stop
        16'd4:
        begin
        state <= stop;
        end

        //load
        16'd5:
        begin
          state <= load;
        end

        //goto
        16'd6:
        begin
          program_counter <= literal_2;
          state <= instruction_fetch;
        end

        //return
        16'd7:
        begin
          program_counter <= operand_a;
          state <= instruction_fetch;
        end

        //add
        16'd8:
        begin
          long_result = operand_a + operand_b;
          result <= long_result[31:0];
          carry[0] <= long_result[32];
          write_enable <= 1;
        end

        //jmp_if_false
        16'd9:
        begin
          if (operand_a == 0) begin
            program_counter <= literal_2;
            state <= instruction_fetch;
          end
        end

        //write
        16'd10:
        begin
          state <= write;
          write_output <= operand_a;
          write_value <= operand_b;
        end

        //read
        16'd11:
        begin
          state <= read;
          read_input <= operand_a;
        end

        //equal
        16'd12:
        begin
          result <= operand_a == operand_b;
          write_enable <= 1;
        end

        //shift_left
        16'd13:
        begin
          if(operand_b < 32) begin
            result <= operand_a << operand_b;
            carry <= operand_a >> (32-operand_b);
          end else begin
            result <= 0;
            carry <= operand_a;
          end
          write_enable <= 1;
        end

        //greater_equal
        16'd14:
        begin
          result <= $signed(operand_a) >= $signed(operand_b);
          write_enable <= 1;
        end

        //jmp_if_true
        16'd15:
        begin
          if (operand_a != 0) begin
            program_counter <= literal_2;
            state <= instruction_fetch;
          end
        end

        //subtract
        16'd16:
        begin
          long_result = operand_a + (~operand_b) + 1;
          result <= long_result[31:0];
          carry[0] <= ~long_result[32];
          write_enable <= 1;
        end

        //unsigned_greater
        16'd17:
        begin
          result <= $unsigned(operand_a) > $unsigned(operand_b);
          write_enable <= 1;
        end

        //unsigned_shift_right
        16'd18:
        begin
          if(operand_b < 32) begin
            result <= operand_a >> operand_b;
            carry <= operand_a << (32-operand_b);
          end else begin
            result <= 0;
            carry <= operand_a;
          end
          write_enable <= 1;
        end

      endcase

    end

    read:
    begin
      case(read_input)
      4:
      begin
        s_input_rs232_rx_ack <= 1;
        if (s_input_rs232_rx_ack && input_rs232_rx_stb) begin
          result <= input_rs232_rx;
          write_enable <= 1;
          s_input_rs232_rx_ack <= 0;
          state <= execute;
        end
      end
      endcase
    end

    write:
    begin
      case(write_output)
      0:
      begin
        s_output_led_r_stb <= 1;
        s_output_led_r <= write_value;
        if (output_led_r_ack && s_output_led_r_stb) begin
          s_output_led_r_stb <= 0;
          state <= execute;
        end
      end
      1:
      begin
        s_output_led_g_stb <= 1;
        s_output_led_g <= write_value;
        if (output_led_g_ack && s_output_led_g_stb) begin
          s_output_led_g_stb <= 0;
          state <= execute;
        end
      end
      2:
      begin
        s_output_led_b_stb <= 1;
        s_output_led_b <= write_value;
        if (output_led_b_ack && s_output_led_b_stb) begin
          s_output_led_b_stb <= 0;
          state <= execute;
        end
      end
      3:
      begin
        s_output_rs232_tx_stb <= 1;
        s_output_rs232_tx <= write_value;
        if (output_rs232_tx_ack && s_output_rs232_tx_stb) begin
          s_output_rs232_tx_stb <= 0;
          state <= execute;
        end
      end
      endcase
    end

    load:
    begin
        result <= load_data;
        write_enable <= 1;
        state <= execute;
    end

    wait_state:
    begin
      if (timer) begin
        timer <= timer - 1;
      end else begin
        state <= execute;
      end
    end

    stop:
    begin
    end

    endcase

    if (rst == 1'b1) begin
      timer <= 0;
      timer_clock <= 0;
      program_counter <= 0;
      address_z_3 <= 0;
      result <= 0;
      a = 0;
      b = 0;
      z = 0;
      state <= instruction_fetch;
      s_input_rs232_rx_ack <= 0;
      s_output_led_r_stb <= 0;
      s_output_led_g_stb <= 0;
      s_output_led_b_stb <= 0;
      s_output_rs232_tx_stb <= 0;
    end
  end
  assign input_rs232_rx_ack = s_input_rs232_rx_ack;
  assign output_led_r_stb = s_output_led_r_stb;
  assign output_led_r = s_output_led_r;
  assign output_led_g_stb = s_output_led_g_stb;
  assign output_led_g = s_output_led_g;
  assign output_led_b_stb = s_output_led_b_stb;
  assign output_led_b = s_output_led_b;
  assign output_rs232_tx_stb = s_output_rs232_tx_stb;
  assign output_rs232_tx = s_output_rs232_tx;

endmodule
