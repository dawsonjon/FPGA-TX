//////////////////////////////////////////////////////////////////////////////
//name : server
//input : input_eth_rx:16
//input : input_socket:16
//output : output_eth_tx:16
//output : output_socket:16
//output : output_rs232_tx:16
//source_file : /media/storage/Projects/Chips-Demo/demo/examples/image_processor/server.c
///======
///
///Created by C2CHIP

module server(input_eth_rx,input_socket,input_eth_rx_stb,input_socket_stb,output_eth_tx_ack,output_socket_ack,output_rs232_tx_ack,clk,rst,output_eth_tx,output_socket,output_rs232_tx,output_eth_tx_stb,output_socket_stb,output_rs232_tx_stb,input_eth_rx_ack,input_socket_ack,exception);
  integer file_count;
  parameter  stop = 3'd0,
  instruction_fetch = 3'd1,
  operand_fetch = 3'd2,
  execute = 3'd3,
  load = 3'd4,
  wait_state = 3'd5,
  read = 3'd6,
  write = 3'd7;
  input [31:0] input_eth_rx;
  input [31:0] input_socket;
  input input_eth_rx_stb;
  input input_socket_stb;
  input output_eth_tx_ack;
  input output_socket_ack;
  input output_rs232_tx_ack;
  input clk;
  input rst;
  output [31:0] output_eth_tx;
  output [31:0] output_socket;
  output [31:0] output_rs232_tx;
  output output_eth_tx_stb;
  output output_socket_stb;
  output output_rs232_tx_stb;
  output input_eth_rx_ack;
  output input_socket_ack;
  reg [15:0] timer;
  reg [15:0] program_counter;
  reg [15:0] program_counter_1;
  reg [15:0] program_counter_2;
  reg [44:0] instruction;
  reg [4:0] opcode_2;
  reg [3:0] a;
  reg [3:0] b;
  reg [3:0] z;
  reg write_enable;
  reg [3:0] address_a_2;
  reg [3:0] address_b_2;
  reg [3:0] address_z_2;
  reg [3:0] address_z_3;
  reg [31:0] load_data;
  reg [31:0] write_output;
  reg [31:0] write_value;
  reg [31:0] read_input;
  reg [31:0] literal_2;
  reg [31:0] a_hi;
  reg [31:0] b_hi;
  reg [31:0] a_lo;
  reg [31:0] b_lo;
  reg [63:0] long_result;
  reg [31:0] result;
  reg [15:0] address;
  reg [31:0] data_out;
  reg [31:0] data_in;
  reg [31:0] carry;
  reg [31:0] s_output_eth_tx_stb;
  reg [31:0] s_output_socket_stb;
  reg [31:0] s_output_rs232_tx_stb;
  reg [31:0] s_output_eth_tx;
  reg [31:0] s_output_socket;
  reg [31:0] s_output_rs232_tx;
  reg [31:0] s_input_eth_rx_ack;
  reg [31:0] s_input_socket_ack;
  reg [7:0] state;
  output reg exception;
  reg [44:0] instructions [5996:0];
  reg [31:0] memory [6143:0];
  reg [31:0] registers [15:0];
  wire [31:0] operand_a;
  wire [31:0] operand_b;
  wire [31:0] register_a;
  wire [31:0] register_b;
  wire [31:0] literal;
  wire [4:0] opcode;
  wire [3:0] address_a;
  wire [3:0] address_b;
  wire [3:0] address_z;
  wire [15:0] load_address;
  wire [15:0] store_address;
  wire [31:0] store_data;
  wire  store_enable;

  //////////////////////////////////////////////////////////////////////////////
  // INSTRUCTION INITIALIZATION                                                 
  //                                                                            
  // Initialise the contents of the instruction memory                          
  //
  // Intruction Set
  // ==============
  // 0 {'literal': True, 'op': 'literal'}
  // 1 {'literal': True, 'op': 'addl'}
  // 2 {'literal': False, 'op': 'store'}
  // 3 {'literal': True, 'op': 'call'}
  // 4 {'literal': False, 'op': 'stop'}
  // 5 {'literal': False, 'op': 'load'}
  // 6 {'literal': True, 'op': 'jmp_if_false'}
  // 7 {'literal': False, 'op': 'equal'}
  // 8 {'literal': True, 'op': 'goto'}
  // 9 {'literal': False, 'op': 'add'}
  // 10 {'literal': False, 'op': 'subtract'}
  // 11 {'literal': False, 'op': 'wait_clocks'}
  // 12 {'literal': False, 'op': 'return'}
  // 13 {'literal': False, 'op': 'write'}
  // 14 {'literal': False, 'op': 'unsigned_shift_right'}
  // 15 {'literal': False, 'op': 'and'}
  // 16 {'literal': False, 'op': 'shift_left'}
  // 17 {'literal': False, 'op': 'or'}
  // 18 {'literal': False, 'op': 'not_equal'}
  // 19 {'literal': False, 'op': 'unsigned_greater_equal'}
  // 20 {'literal': False, 'op': 'unsigned_greater'}
  // 21 {'literal': False, 'op': 'ready'}
  // 22 {'literal': False, 'op': 'read'}
  // 23 {'literal': False, 'op': 'int_to_long'}
  // 24 {'literal': False, 'op': 'add_with_carry'}
  // 25 {'literal': False, 'op': 'not'}
  // 26 {'literal': False, 'op': 'output_ready'}
  // 27 {'literal': True, 'op': 'jmp_if_true'}
  // Intructions
  // ===========
  
  initial
  begin
    instructions[0] = {5'd0, 4'd3, 4'd0, 32'd0};//{'literal': 0, 'z': 3, 'op': 'literal'}
    instructions[1] = {5'd0, 4'd4, 4'd0, 32'd0};//{'literal': 0, 'z': 4, 'op': 'literal'}
    instructions[2] = {5'd1, 4'd3, 4'd3, 32'd2744};//{'a': 3, 'literal': 2744, 'z': 3, 'op': 'addl'}
    instructions[3] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[4] = {5'd0, 4'd2, 4'd0, 32'd1};//{'literal': 1, 'z': 2, 'op': 'literal'}
    instructions[5] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[6] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[7] = {5'd0, 4'd2, 4'd0, 32'd2};//{'literal': 2, 'z': 2, 'op': 'literal'}
    instructions[8] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[9] = {5'd0, 4'd8, 4'd0, 32'd69};//{'literal': 69, 'z': 8, 'op': 'literal'}
    instructions[10] = {5'd0, 4'd2, 4'd0, 32'd3};//{'literal': 3, 'z': 2, 'op': 'literal'}
    instructions[11] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[12] = {5'd0, 4'd8, 4'd0, 32'd83};//{'literal': 83, 'z': 8, 'op': 'literal'}
    instructions[13] = {5'd0, 4'd2, 4'd0, 32'd4};//{'literal': 4, 'z': 2, 'op': 'literal'}
    instructions[14] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[15] = {5'd0, 4'd8, 4'd0, 32'd84};//{'literal': 84, 'z': 8, 'op': 'literal'}
    instructions[16] = {5'd0, 4'd2, 4'd0, 32'd5};//{'literal': 5, 'z': 2, 'op': 'literal'}
    instructions[17] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[18] = {5'd0, 4'd8, 4'd0, 32'd65};//{'literal': 65, 'z': 8, 'op': 'literal'}
    instructions[19] = {5'd0, 4'd2, 4'd0, 32'd6};//{'literal': 6, 'z': 2, 'op': 'literal'}
    instructions[20] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[21] = {5'd0, 4'd8, 4'd0, 32'd66};//{'literal': 66, 'z': 8, 'op': 'literal'}
    instructions[22] = {5'd0, 4'd2, 4'd0, 32'd7};//{'literal': 7, 'z': 2, 'op': 'literal'}
    instructions[23] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[24] = {5'd0, 4'd8, 4'd0, 32'd76};//{'literal': 76, 'z': 8, 'op': 'literal'}
    instructions[25] = {5'd0, 4'd2, 4'd0, 32'd8};//{'literal': 8, 'z': 2, 'op': 'literal'}
    instructions[26] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[27] = {5'd0, 4'd8, 4'd0, 32'd73};//{'literal': 73, 'z': 8, 'op': 'literal'}
    instructions[28] = {5'd0, 4'd2, 4'd0, 32'd9};//{'literal': 9, 'z': 2, 'op': 'literal'}
    instructions[29] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[30] = {5'd0, 4'd8, 4'd0, 32'd83};//{'literal': 83, 'z': 8, 'op': 'literal'}
    instructions[31] = {5'd0, 4'd2, 4'd0, 32'd10};//{'literal': 10, 'z': 2, 'op': 'literal'}
    instructions[32] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[33] = {5'd0, 4'd8, 4'd0, 32'd72};//{'literal': 72, 'z': 8, 'op': 'literal'}
    instructions[34] = {5'd0, 4'd2, 4'd0, 32'd11};//{'literal': 11, 'z': 2, 'op': 'literal'}
    instructions[35] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[36] = {5'd0, 4'd8, 4'd0, 32'd69};//{'literal': 69, 'z': 8, 'op': 'literal'}
    instructions[37] = {5'd0, 4'd2, 4'd0, 32'd12};//{'literal': 12, 'z': 2, 'op': 'literal'}
    instructions[38] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[39] = {5'd0, 4'd8, 4'd0, 32'd68};//{'literal': 68, 'z': 8, 'op': 'literal'}
    instructions[40] = {5'd0, 4'd2, 4'd0, 32'd13};//{'literal': 13, 'z': 2, 'op': 'literal'}
    instructions[41] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[42] = {5'd0, 4'd8, 4'd0, 32'd10};//{'literal': 10, 'z': 8, 'op': 'literal'}
    instructions[43] = {5'd0, 4'd2, 4'd0, 32'd14};//{'literal': 14, 'z': 2, 'op': 'literal'}
    instructions[44] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[45] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[46] = {5'd0, 4'd2, 4'd0, 32'd15};//{'literal': 15, 'z': 2, 'op': 'literal'}
    instructions[47] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[48] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[49] = {5'd0, 4'd2, 4'd0, 32'd16};//{'literal': 16, 'z': 2, 'op': 'literal'}
    instructions[50] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[51] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[52] = {5'd0, 4'd2, 4'd0, 32'd33};//{'literal': 33, 'z': 2, 'op': 'literal'}
    instructions[53] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[54] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[55] = {5'd0, 4'd2, 4'd0, 32'd34};//{'literal': 34, 'z': 2, 'op': 'literal'}
    instructions[56] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[57] = {5'd0, 4'd8, 4'd0, 32'd80};//{'literal': 80, 'z': 8, 'op': 'literal'}
    instructions[58] = {5'd0, 4'd2, 4'd0, 32'd35};//{'literal': 35, 'z': 2, 'op': 'literal'}
    instructions[59] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[60] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[61] = {5'd0, 4'd2, 4'd0, 32'd36};//{'literal': 36, 'z': 2, 'op': 'literal'}
    instructions[62] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[63] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[64] = {5'd0, 4'd2, 4'd0, 32'd37};//{'literal': 37, 'z': 2, 'op': 'literal'}
    instructions[65] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[66] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[67] = {5'd0, 4'd9, 4'd0, 32'd0};//{'literal': 0, 'z': 9, 'op': 'literal'}
    instructions[68] = {5'd0, 4'd2, 4'd0, 32'd38};//{'literal': 38, 'z': 2, 'op': 'literal'}
    instructions[69] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[70] = {5'd1, 4'd2, 4'd2, 32'd1};//{'a': 2, 'literal': 1, 'z': 2, 'op': 'addl'}
    instructions[71] = {5'd2, 4'd0, 4'd2, 32'd9};//{'a': 2, 'b': 9, 'op': 'store'}
    instructions[72] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[73] = {5'd0, 4'd2, 4'd0, 32'd40};//{'literal': 40, 'z': 2, 'op': 'literal'}
    instructions[74] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[75] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[76] = {5'd0, 4'd2, 4'd0, 32'd41};//{'literal': 41, 'z': 2, 'op': 'literal'}
    instructions[77] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[78] = {5'd0, 4'd8, 4'd0, 32'd49320};//{'literal': 49320, 'z': 8, 'op': 'literal'}
    instructions[79] = {5'd0, 4'd2, 4'd0, 32'd44};//{'literal': 44, 'z': 2, 'op': 'literal'}
    instructions[80] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[81] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[82] = {5'd0, 4'd2, 4'd0, 32'd45};//{'literal': 45, 'z': 2, 'op': 'literal'}
    instructions[83] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[84] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[85] = {5'd0, 4'd2, 4'd0, 32'd46};//{'literal': 46, 'z': 2, 'op': 'literal'}
    instructions[86] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[87] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[88] = {5'd0, 4'd2, 4'd0, 32'd47};//{'literal': 47, 'z': 2, 'op': 'literal'}
    instructions[89] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[90] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[91] = {5'd0, 4'd2, 4'd0, 32'd48};//{'literal': 48, 'z': 2, 'op': 'literal'}
    instructions[92] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[93] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[94] = {5'd0, 4'd2, 4'd0, 32'd49};//{'literal': 49, 'z': 2, 'op': 'literal'}
    instructions[95] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[96] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[97] = {5'd0, 4'd2, 4'd0, 32'd50};//{'literal': 50, 'z': 2, 'op': 'literal'}
    instructions[98] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[99] = {5'd0, 4'd8, 4'd0, 32'd1024};//{'literal': 1024, 'z': 8, 'op': 'literal'}
    instructions[100] = {5'd0, 4'd2, 4'd0, 32'd51};//{'literal': 51, 'z': 2, 'op': 'literal'}
    instructions[101] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[102] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[103] = {5'd0, 4'd2, 4'd0, 32'd52};//{'literal': 52, 'z': 2, 'op': 'literal'}
    instructions[104] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[105] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[106] = {5'd0, 4'd2, 4'd0, 32'd53};//{'literal': 53, 'z': 2, 'op': 'literal'}
    instructions[107] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[108] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[109] = {5'd0, 4'd2, 4'd0, 32'd1078};//{'literal': 1078, 'z': 2, 'op': 'literal'}
    instructions[110] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[111] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[112] = {5'd0, 4'd2, 4'd0, 32'd1079};//{'literal': 1079, 'z': 2, 'op': 'literal'}
    instructions[113] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[114] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[115] = {5'd0, 4'd2, 4'd0, 32'd1080};//{'literal': 1080, 'z': 2, 'op': 'literal'}
    instructions[116] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[117] = {5'd0, 4'd8, 4'd0, 32'd76};//{'literal': 76, 'z': 8, 'op': 'literal'}
    instructions[118] = {5'd0, 4'd2, 4'd0, 32'd1082};//{'literal': 1082, 'z': 2, 'op': 'literal'}
    instructions[119] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[120] = {5'd0, 4'd8, 4'd0, 32'd73};//{'literal': 73, 'z': 8, 'op': 'literal'}
    instructions[121] = {5'd0, 4'd2, 4'd0, 32'd1083};//{'literal': 1083, 'z': 2, 'op': 'literal'}
    instructions[122] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[123] = {5'd0, 4'd8, 4'd0, 32'd83};//{'literal': 83, 'z': 8, 'op': 'literal'}
    instructions[124] = {5'd0, 4'd2, 4'd0, 32'd1084};//{'literal': 1084, 'z': 2, 'op': 'literal'}
    instructions[125] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[126] = {5'd0, 4'd8, 4'd0, 32'd84};//{'literal': 84, 'z': 8, 'op': 'literal'}
    instructions[127] = {5'd0, 4'd2, 4'd0, 32'd1085};//{'literal': 1085, 'z': 2, 'op': 'literal'}
    instructions[128] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[129] = {5'd0, 4'd8, 4'd0, 32'd69};//{'literal': 69, 'z': 8, 'op': 'literal'}
    instructions[130] = {5'd0, 4'd2, 4'd0, 32'd1086};//{'literal': 1086, 'z': 2, 'op': 'literal'}
    instructions[131] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[132] = {5'd0, 4'd8, 4'd0, 32'd78};//{'literal': 78, 'z': 8, 'op': 'literal'}
    instructions[133] = {5'd0, 4'd2, 4'd0, 32'd1087};//{'literal': 1087, 'z': 2, 'op': 'literal'}
    instructions[134] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[135] = {5'd0, 4'd8, 4'd0, 32'd10};//{'literal': 10, 'z': 8, 'op': 'literal'}
    instructions[136] = {5'd0, 4'd2, 4'd0, 32'd1088};//{'literal': 1088, 'z': 2, 'op': 'literal'}
    instructions[137] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[138] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[139] = {5'd0, 4'd2, 4'd0, 32'd1089};//{'literal': 1089, 'z': 2, 'op': 'literal'}
    instructions[140] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[141] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[142] = {5'd0, 4'd2, 4'd0, 32'd1090};//{'literal': 1090, 'z': 2, 'op': 'literal'}
    instructions[143] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[144] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[145] = {5'd0, 4'd2, 4'd0, 32'd1091};//{'literal': 1091, 'z': 2, 'op': 'literal'}
    instructions[146] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[147] = {5'd0, 4'd8, 4'd0, 32'd515};//{'literal': 515, 'z': 8, 'op': 'literal'}
    instructions[148] = {5'd0, 4'd2, 4'd0, 32'd1109};//{'literal': 1109, 'z': 2, 'op': 'literal'}
    instructions[149] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[150] = {5'd0, 4'd8, 4'd0, 32'd87};//{'literal': 87, 'z': 8, 'op': 'literal'}
    instructions[151] = {5'd0, 4'd2, 4'd0, 32'd1110};//{'literal': 1110, 'z': 2, 'op': 'literal'}
    instructions[152] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[153] = {5'd0, 4'd8, 4'd0, 32'd65};//{'literal': 65, 'z': 8, 'op': 'literal'}
    instructions[154] = {5'd0, 4'd2, 4'd0, 32'd1111};//{'literal': 1111, 'z': 2, 'op': 'literal'}
    instructions[155] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[156] = {5'd0, 4'd8, 4'd0, 32'd73};//{'literal': 73, 'z': 8, 'op': 'literal'}
    instructions[157] = {5'd0, 4'd2, 4'd0, 32'd1112};//{'literal': 1112, 'z': 2, 'op': 'literal'}
    instructions[158] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[159] = {5'd0, 4'd8, 4'd0, 32'd84};//{'literal': 84, 'z': 8, 'op': 'literal'}
    instructions[160] = {5'd0, 4'd2, 4'd0, 32'd1113};//{'literal': 1113, 'z': 2, 'op': 'literal'}
    instructions[161] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[162] = {5'd0, 4'd8, 4'd0, 32'd32};//{'literal': 32, 'z': 8, 'op': 'literal'}
    instructions[163] = {5'd0, 4'd2, 4'd0, 32'd1114};//{'literal': 1114, 'z': 2, 'op': 'literal'}
    instructions[164] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[165] = {5'd0, 4'd8, 4'd0, 32'd67};//{'literal': 67, 'z': 8, 'op': 'literal'}
    instructions[166] = {5'd0, 4'd2, 4'd0, 32'd1115};//{'literal': 1115, 'z': 2, 'op': 'literal'}
    instructions[167] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[168] = {5'd0, 4'd8, 4'd0, 32'd76};//{'literal': 76, 'z': 8, 'op': 'literal'}
    instructions[169] = {5'd0, 4'd2, 4'd0, 32'd1116};//{'literal': 1116, 'z': 2, 'op': 'literal'}
    instructions[170] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[171] = {5'd0, 4'd8, 4'd0, 32'd79};//{'literal': 79, 'z': 8, 'op': 'literal'}
    instructions[172] = {5'd0, 4'd2, 4'd0, 32'd1117};//{'literal': 1117, 'z': 2, 'op': 'literal'}
    instructions[173] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[174] = {5'd0, 4'd8, 4'd0, 32'd83};//{'literal': 83, 'z': 8, 'op': 'literal'}
    instructions[175] = {5'd0, 4'd2, 4'd0, 32'd1118};//{'literal': 1118, 'z': 2, 'op': 'literal'}
    instructions[176] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[177] = {5'd0, 4'd8, 4'd0, 32'd69};//{'literal': 69, 'z': 8, 'op': 'literal'}
    instructions[178] = {5'd0, 4'd2, 4'd0, 32'd1119};//{'literal': 1119, 'z': 2, 'op': 'literal'}
    instructions[179] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[180] = {5'd0, 4'd8, 4'd0, 32'd10};//{'literal': 10, 'z': 8, 'op': 'literal'}
    instructions[181] = {5'd0, 4'd2, 4'd0, 32'd1120};//{'literal': 1120, 'z': 2, 'op': 'literal'}
    instructions[182] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[183] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[184] = {5'd0, 4'd2, 4'd0, 32'd1121};//{'literal': 1121, 'z': 2, 'op': 'literal'}
    instructions[185] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[186] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[187] = {5'd0, 4'd2, 4'd0, 32'd1122};//{'literal': 1122, 'z': 2, 'op': 'literal'}
    instructions[188] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[189] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[190] = {5'd0, 4'd2, 4'd0, 32'd1123};//{'literal': 1123, 'z': 2, 'op': 'literal'}
    instructions[191] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[192] = {5'd0, 4'd8, 4'd0, 32'd257};//{'literal': 257, 'z': 8, 'op': 'literal'}
    instructions[193] = {5'd0, 4'd2, 4'd0, 32'd1124};//{'literal': 1124, 'z': 2, 'op': 'literal'}
    instructions[194] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[195] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[196] = {5'd0, 4'd2, 4'd0, 32'd1125};//{'literal': 1125, 'z': 2, 'op': 'literal'}
    instructions[197] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[198] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[199] = {5'd0, 4'd2, 4'd0, 32'd1126};//{'literal': 1126, 'z': 2, 'op': 'literal'}
    instructions[200] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[201] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[202] = {5'd0, 4'd2, 4'd0, 32'd1127};//{'literal': 1127, 'z': 2, 'op': 'literal'}
    instructions[203] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[204] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[205] = {5'd0, 4'd2, 4'd0, 32'd1128};//{'literal': 1128, 'z': 2, 'op': 'literal'}
    instructions[206] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[207] = {5'd0, 4'd8, 4'd0, 32'd4};//{'literal': 4, 'z': 8, 'op': 'literal'}
    instructions[208] = {5'd0, 4'd2, 4'd0, 32'd1129};//{'literal': 1129, 'z': 2, 'op': 'literal'}
    instructions[209] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[210] = {5'd0, 4'd8, 4'd0, 32'd3};//{'literal': 3, 'z': 8, 'op': 'literal'}
    instructions[211] = {5'd0, 4'd2, 4'd0, 32'd2154};//{'literal': 2154, 'z': 2, 'op': 'literal'}
    instructions[212] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[213] = {5'd0, 4'd8, 4'd0, 32'd83};//{'literal': 83, 'z': 8, 'op': 'literal'}
    instructions[214] = {5'd0, 4'd2, 4'd0, 32'd2685};//{'literal': 2685, 'z': 2, 'op': 'literal'}
    instructions[215] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[216] = {5'd0, 4'd8, 4'd0, 32'd89};//{'literal': 89, 'z': 8, 'op': 'literal'}
    instructions[217] = {5'd0, 4'd2, 4'd0, 32'd2686};//{'literal': 2686, 'z': 2, 'op': 'literal'}
    instructions[218] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[219] = {5'd0, 4'd8, 4'd0, 32'd78};//{'literal': 78, 'z': 8, 'op': 'literal'}
    instructions[220] = {5'd0, 4'd2, 4'd0, 32'd2687};//{'literal': 2687, 'z': 2, 'op': 'literal'}
    instructions[221] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[222] = {5'd0, 4'd8, 4'd0, 32'd32};//{'literal': 32, 'z': 8, 'op': 'literal'}
    instructions[223] = {5'd0, 4'd2, 4'd0, 32'd2688};//{'literal': 2688, 'z': 2, 'op': 'literal'}
    instructions[224] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[225] = {5'd0, 4'd8, 4'd0, 32'd82};//{'literal': 82, 'z': 8, 'op': 'literal'}
    instructions[226] = {5'd0, 4'd2, 4'd0, 32'd2689};//{'literal': 2689, 'z': 2, 'op': 'literal'}
    instructions[227] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[228] = {5'd0, 4'd8, 4'd0, 32'd69};//{'literal': 69, 'z': 8, 'op': 'literal'}
    instructions[229] = {5'd0, 4'd2, 4'd0, 32'd2690};//{'literal': 2690, 'z': 2, 'op': 'literal'}
    instructions[230] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[231] = {5'd0, 4'd8, 4'd0, 32'd67};//{'literal': 67, 'z': 8, 'op': 'literal'}
    instructions[232] = {5'd0, 4'd2, 4'd0, 32'd2691};//{'literal': 2691, 'z': 2, 'op': 'literal'}
    instructions[233] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[234] = {5'd0, 4'd8, 4'd0, 32'd69};//{'literal': 69, 'z': 8, 'op': 'literal'}
    instructions[235] = {5'd0, 4'd2, 4'd0, 32'd2692};//{'literal': 2692, 'z': 2, 'op': 'literal'}
    instructions[236] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[237] = {5'd0, 4'd8, 4'd0, 32'd73};//{'literal': 73, 'z': 8, 'op': 'literal'}
    instructions[238] = {5'd0, 4'd2, 4'd0, 32'd2693};//{'literal': 2693, 'z': 2, 'op': 'literal'}
    instructions[239] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[240] = {5'd0, 4'd8, 4'd0, 32'd86};//{'literal': 86, 'z': 8, 'op': 'literal'}
    instructions[241] = {5'd0, 4'd2, 4'd0, 32'd2694};//{'literal': 2694, 'z': 2, 'op': 'literal'}
    instructions[242] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[243] = {5'd0, 4'd8, 4'd0, 32'd69};//{'literal': 69, 'z': 8, 'op': 'literal'}
    instructions[244] = {5'd0, 4'd2, 4'd0, 32'd2695};//{'literal': 2695, 'z': 2, 'op': 'literal'}
    instructions[245] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[246] = {5'd0, 4'd8, 4'd0, 32'd68};//{'literal': 68, 'z': 8, 'op': 'literal'}
    instructions[247] = {5'd0, 4'd2, 4'd0, 32'd2696};//{'literal': 2696, 'z': 2, 'op': 'literal'}
    instructions[248] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[249] = {5'd0, 4'd8, 4'd0, 32'd10};//{'literal': 10, 'z': 8, 'op': 'literal'}
    instructions[250] = {5'd0, 4'd2, 4'd0, 32'd2697};//{'literal': 2697, 'z': 2, 'op': 'literal'}
    instructions[251] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[252] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[253] = {5'd0, 4'd2, 4'd0, 32'd2698};//{'literal': 2698, 'z': 2, 'op': 'literal'}
    instructions[254] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[255] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[256] = {5'd0, 4'd2, 4'd0, 32'd2699};//{'literal': 2699, 'z': 2, 'op': 'literal'}
    instructions[257] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[258] = {5'd0, 4'd8, 4'd0, 32'd1029};//{'literal': 1029, 'z': 8, 'op': 'literal'}
    instructions[259] = {5'd0, 4'd2, 4'd0, 32'd2702};//{'literal': 2702, 'z': 2, 'op': 'literal'}
    instructions[260] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[261] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[262] = {5'd0, 4'd2, 4'd0, 32'd2703};//{'literal': 2703, 'z': 2, 'op': 'literal'}
    instructions[263] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[264] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[265] = {5'd0, 4'd2, 4'd0, 32'd2704};//{'literal': 2704, 'z': 2, 'op': 'literal'}
    instructions[266] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[267] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[268] = {5'd0, 4'd2, 4'd0, 32'd2721};//{'literal': 2721, 'z': 2, 'op': 'literal'}
    instructions[269] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[270] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[271] = {5'd0, 4'd2, 4'd0, 32'd2722};//{'literal': 2722, 'z': 2, 'op': 'literal'}
    instructions[272] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[273] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[274] = {5'd0, 4'd2, 4'd0, 32'd2723};//{'literal': 2723, 'z': 2, 'op': 'literal'}
    instructions[275] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[276] = {5'd0, 4'd8, 4'd0, 32'd1024};//{'literal': 1024, 'z': 8, 'op': 'literal'}
    instructions[277] = {5'd0, 4'd2, 4'd0, 32'd2724};//{'literal': 2724, 'z': 2, 'op': 'literal'}
    instructions[278] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[279] = {5'd0, 4'd8, 4'd0, 32'd2};//{'literal': 2, 'z': 8, 'op': 'literal'}
    instructions[280] = {5'd0, 4'd2, 4'd0, 32'd2725};//{'literal': 2725, 'z': 2, 'op': 'literal'}
    instructions[281] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[282] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[283] = {5'd0, 4'd2, 4'd0, 32'd2726};//{'literal': 2726, 'z': 2, 'op': 'literal'}
    instructions[284] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[285] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[286] = {5'd0, 4'd2, 4'd0, 32'd2727};//{'literal': 2727, 'z': 2, 'op': 'literal'}
    instructions[287] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[288] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[289] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[290] = {5'd3, 4'd6, 4'd0, 32'd292};//{'z': 6, 'label': 292, 'op': 'call'}
    instructions[291] = {5'd4, 4'd0, 4'd0, 32'd0};//{'op': 'stop'}
    instructions[292] = {5'd1, 4'd3, 4'd3, 32'd2102};//{'a': 3, 'literal': 2102, 'z': 3, 'op': 'addl'}
    instructions[293] = {5'd0, 4'd8, 4'd0, 32'd27};//{'literal': 27, 'z': 8, 'op': 'literal'}
    instructions[294] = {5'd1, 4'd2, 4'd4, 32'd2048};//{'a': 4, 'literal': 2048, 'z': 2, 'op': 'addl'}
    instructions[295] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[296] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[297] = {5'd1, 4'd2, 4'd4, 32'd2049};//{'a': 4, 'literal': 2049, 'z': 2, 'op': 'addl'}
    instructions[298] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[299] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[300] = {5'd1, 4'd2, 4'd4, 32'd2050};//{'a': 4, 'literal': 2050, 'z': 2, 'op': 'addl'}
    instructions[301] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[302] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[303] = {5'd1, 4'd2, 4'd4, 32'd2051};//{'a': 4, 'literal': 2051, 'z': 2, 'op': 'addl'}
    instructions[304] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[305] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[306] = {5'd1, 4'd2, 4'd4, 32'd2052};//{'a': 4, 'literal': 2052, 'z': 2, 'op': 'addl'}
    instructions[307] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[308] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[309] = {5'd1, 4'd2, 4'd4, 32'd2053};//{'a': 4, 'literal': 2053, 'z': 2, 'op': 'addl'}
    instructions[310] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[311] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[312] = {5'd1, 4'd2, 4'd4, 32'd2054};//{'a': 4, 'literal': 2054, 'z': 2, 'op': 'addl'}
    instructions[313] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[314] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[315] = {5'd0, 4'd2, 4'd0, 32'd2703};//{'literal': 2703, 'z': 2, 'op': 'literal'}
    instructions[316] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[317] = {5'd0, 4'd8, 4'd0, 32'd1129};//{'literal': 1129, 'z': 8, 'op': 'literal'}
    instructions[318] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[319] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[320] = {5'd0, 4'd2, 4'd0, 32'd47};//{'literal': 47, 'z': 2, 'op': 'literal'}
    instructions[321] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[322] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[323] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[324] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[325] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[326] = {5'd0, 4'd8, 4'd0, 32'd1082};//{'literal': 1082, 'z': 8, 'op': 'literal'}
    instructions[327] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[328] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[329] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[330] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[331] = {5'd3, 4'd6, 4'd0, 32'd1264};//{'z': 6, 'label': 1264, 'op': 'call'}
    instructions[332] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[333] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[334] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[335] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[336] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[337] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[338] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[339] = {5'd0, 4'd2, 4'd0, 32'd41};//{'literal': 41, 'z': 2, 'op': 'literal'}
    instructions[340] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[341] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[342] = {5'd0, 4'd2, 4'd0, 32'd1079};//{'literal': 1079, 'z': 2, 'op': 'literal'}
    instructions[343] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[344] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[345] = {5'd0, 4'd2, 4'd0, 32'd2704};//{'literal': 2704, 'z': 2, 'op': 'literal'}
    instructions[346] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[347] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[348] = {5'd0, 4'd2, 4'd0, 32'd2699};//{'literal': 2699, 'z': 2, 'op': 'literal'}
    instructions[349] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[350] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[351] = {5'd0, 4'd2, 4'd0, 32'd34};//{'literal': 34, 'z': 2, 'op': 'literal'}
    instructions[352] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[353] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[354] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[355] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[356] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[357] = {5'd1, 4'd8, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 8, 'op': 'addl'}
    instructions[358] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[359] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[360] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[361] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[362] = {5'd3, 4'd6, 4'd0, 32'd1352};//{'z': 6, 'label': 1352, 'op': 'call'}
    instructions[363] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[364] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[365] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[366] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[367] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[368] = {5'd0, 4'd2, 4'd0, 32'd2701};//{'literal': 2701, 'z': 2, 'op': 'literal'}
    instructions[369] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[370] = {5'd1, 4'd2, 4'd4, 32'd2051};//{'a': 4, 'literal': 2051, 'z': 2, 'op': 'addl'}
    instructions[371] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[372] = {5'd1, 4'd8, 4'd4, 32'd2051};//{'a': 4, 'literal': 2051, 'z': 8, 'op': 'addl'}
    instructions[373] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[374] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[375] = {5'd6, 4'd0, 4'd8, 32'd385};//{'a': 8, 'label': 385, 'op': 'jmp_if_false'}
    instructions[376] = {5'd0, 4'd8, 4'd0, 32'd80};//{'literal': 80, 'z': 8, 'op': 'literal'}
    instructions[377] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[378] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[379] = {5'd0, 4'd8, 4'd0, 32'd2726};//{'literal': 2726, 'z': 8, 'op': 'literal'}
    instructions[380] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[381] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[382] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[383] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[384] = {5'd7, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'equal'}
    instructions[385] = {5'd6, 4'd0, 4'd8, 32'd389};//{'a': 8, 'label': 389, 'op': 'jmp_if_false'}
    instructions[386] = {5'd0, 4'd8, 4'd0, 32'd1128};//{'literal': 1128, 'z': 8, 'op': 'literal'}
    instructions[387] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[388] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[389] = {5'd6, 4'd0, 4'd8, 32'd392};//{'a': 8, 'label': 392, 'op': 'jmp_if_false'}
    instructions[390] = {5'd8, 4'd0, 4'd0, 32'd393};//{'label': 393, 'op': 'goto'}
    instructions[391] = {5'd8, 4'd0, 4'd0, 32'd392};//{'label': 392, 'op': 'goto'}
    instructions[392] = {5'd8, 4'd0, 4'd0, 32'd353};//{'label': 353, 'op': 'goto'}
    instructions[393] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[394] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[395] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[396] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[397] = {5'd0, 4'd8, 4'd0, 32'd2685};//{'literal': 2685, 'z': 8, 'op': 'literal'}
    instructions[398] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[399] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[400] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[401] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[402] = {5'd3, 4'd6, 4'd0, 32'd1264};//{'z': 6, 'label': 1264, 'op': 'call'}
    instructions[403] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[404] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[405] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[406] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[407] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[408] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[409] = {5'd1, 4'd8, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 8, 'op': 'addl'}
    instructions[410] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[411] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[412] = {5'd0, 4'd8, 4'd0, 32'd13};//{'literal': 13, 'z': 8, 'op': 'literal'}
    instructions[413] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[414] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[415] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[416] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[417] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[418] = {5'd0, 4'd2, 4'd0, 32'd45};//{'literal': 45, 'z': 2, 'op': 'literal'}
    instructions[419] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[420] = {5'd1, 4'd8, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 8, 'op': 'addl'}
    instructions[421] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[422] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[423] = {5'd0, 4'd8, 4'd0, 32'd14};//{'literal': 14, 'z': 8, 'op': 'literal'}
    instructions[424] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[425] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[426] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[427] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[428] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[429] = {5'd0, 4'd2, 4'd0, 32'd1126};//{'literal': 1126, 'z': 2, 'op': 'literal'}
    instructions[430] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[431] = {5'd0, 4'd8, 4'd0, 32'd40};//{'literal': 40, 'z': 8, 'op': 'literal'}
    instructions[432] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[433] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[434] = {5'd0, 4'd2, 4'd0, 32'd1078};//{'literal': 1078, 'z': 2, 'op': 'literal'}
    instructions[435] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[436] = {5'd0, 4'd8, 4'd0, 32'd80};//{'literal': 80, 'z': 8, 'op': 'literal'}
    instructions[437] = {5'd0, 4'd2, 4'd0, 32'd1091};//{'literal': 1091, 'z': 2, 'op': 'literal'}
    instructions[438] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[439] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[440] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[441] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[442] = {5'd0, 4'd8, 4'd0, 32'd2};//{'literal': 2, 'z': 8, 'op': 'literal'}
    instructions[443] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[444] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[445] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[446] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[447] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[448] = {5'd0, 4'd2, 4'd0, 32'd46};//{'literal': 46, 'z': 2, 'op': 'literal'}
    instructions[449] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[450] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[451] = {5'd0, 4'd2, 4'd0, 32'd1079};//{'literal': 1079, 'z': 2, 'op': 'literal'}
    instructions[452] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[453] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[454] = {5'd0, 4'd2, 4'd0, 32'd2699};//{'literal': 2699, 'z': 2, 'op': 'literal'}
    instructions[455] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[456] = {5'd0, 4'd8, 4'd0, 32'd10000};//{'literal': 10000, 'z': 8, 'op': 'literal'}
    instructions[457] = {5'd1, 4'd2, 4'd4, 32'd2050};//{'a': 4, 'literal': 2050, 'z': 2, 'op': 'addl'}
    instructions[458] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[459] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[460] = {5'd1, 4'd2, 4'd4, 32'd2052};//{'a': 4, 'literal': 2052, 'z': 2, 'op': 'addl'}
    instructions[461] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[462] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[463] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[464] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[465] = {5'd1, 4'd8, 4'd4, 32'd2052};//{'a': 4, 'literal': 2052, 'z': 8, 'op': 'addl'}
    instructions[466] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[467] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[468] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[469] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[470] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[471] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[472] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[473] = {5'd1, 4'd8, 4'd4, 32'd2052};//{'a': 4, 'literal': 2052, 'z': 8, 'op': 'addl'}
    instructions[474] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[475] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[476] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[477] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[478] = {5'd10, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'subtract'}
    instructions[479] = {5'd1, 4'd2, 4'd4, 32'd2052};//{'a': 4, 'literal': 2052, 'z': 2, 'op': 'addl'}
    instructions[480] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[481] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[482] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[483] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[484] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[485] = {5'd7, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'equal'}
    instructions[486] = {5'd6, 4'd0, 4'd8, 32'd537};//{'a': 8, 'label': 537, 'op': 'jmp_if_false'}
    instructions[487] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[488] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[489] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[490] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[491] = {5'd1, 4'd8, 4'd4, 32'd1024};//{'a': 4, 'literal': 1024, 'z': 8, 'op': 'addl'}
    instructions[492] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[493] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[494] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[495] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[496] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[497] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[498] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[499] = {5'd3, 4'd6, 4'd0, 32'd4384};//{'z': 6, 'label': 4384, 'op': 'call'}
    instructions[500] = {5'd1, 4'd3, 4'd3, -32'd2};//{'a': 3, 'literal': -2, 'z': 3, 'op': 'addl'}
    instructions[501] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[502] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[503] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[504] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[505] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[506] = {5'd0, 4'd8, 4'd0, 32'd10};//{'literal': 10, 'z': 8, 'op': 'literal'}
    instructions[507] = {5'd1, 4'd2, 4'd4, 32'd2052};//{'a': 4, 'literal': 2052, 'z': 2, 'op': 'addl'}
    instructions[508] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[509] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[510] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[511] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[512] = {5'd1, 4'd8, 4'd4, 32'd2050};//{'a': 4, 'literal': 2050, 'z': 8, 'op': 'addl'}
    instructions[513] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[514] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[515] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[516] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[517] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[518] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[519] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[520] = {5'd1, 4'd8, 4'd4, 32'd2050};//{'a': 4, 'literal': 2050, 'z': 8, 'op': 'addl'}
    instructions[521] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[522] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[523] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[524] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[525] = {5'd10, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'subtract'}
    instructions[526] = {5'd1, 4'd2, 4'd4, 32'd2050};//{'a': 4, 'literal': 2050, 'z': 2, 'op': 'addl'}
    instructions[527] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[528] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[529] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[530] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[531] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[532] = {5'd7, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'equal'}
    instructions[533] = {5'd6, 4'd0, 4'd8, 32'd536};//{'a': 8, 'label': 536, 'op': 'jmp_if_false'}
    instructions[534] = {5'd8, 4'd0, 4'd0, 32'd589};//{'label': 589, 'op': 'goto'}
    instructions[535] = {5'd8, 4'd0, 4'd0, 32'd536};//{'label': 536, 'op': 'goto'}
    instructions[536] = {5'd8, 4'd0, 4'd0, 32'd537};//{'label': 537, 'op': 'goto'}
    instructions[537] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[538] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[539] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[540] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[541] = {5'd1, 4'd8, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 8, 'op': 'addl'}
    instructions[542] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[543] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[544] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[545] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[546] = {5'd3, 4'd6, 4'd0, 32'd1352};//{'z': 6, 'label': 1352, 'op': 'call'}
    instructions[547] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[548] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[549] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[550] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[551] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[552] = {5'd0, 4'd2, 4'd0, 32'd2701};//{'literal': 2701, 'z': 2, 'op': 'literal'}
    instructions[553] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[554] = {5'd1, 4'd2, 4'd4, 32'd2051};//{'a': 4, 'literal': 2051, 'z': 2, 'op': 'addl'}
    instructions[555] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[556] = {5'd1, 4'd8, 4'd4, 32'd2051};//{'a': 4, 'literal': 2051, 'z': 8, 'op': 'addl'}
    instructions[557] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[558] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[559] = {5'd6, 4'd0, 4'd8, 32'd569};//{'a': 8, 'label': 569, 'op': 'jmp_if_false'}
    instructions[560] = {5'd0, 4'd8, 4'd0, 32'd80};//{'literal': 80, 'z': 8, 'op': 'literal'}
    instructions[561] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[562] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[563] = {5'd0, 4'd8, 4'd0, 32'd2726};//{'literal': 2726, 'z': 8, 'op': 'literal'}
    instructions[564] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[565] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[566] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[567] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[568] = {5'd7, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'equal'}
    instructions[569] = {5'd6, 4'd0, 4'd8, 32'd581};//{'a': 8, 'label': 581, 'op': 'jmp_if_false'}
    instructions[570] = {5'd0, 4'd8, 4'd0, 32'd1078};//{'literal': 1078, 'z': 8, 'op': 'literal'}
    instructions[571] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[572] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[573] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[574] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[575] = {5'd0, 4'd8, 4'd0, 32'd40};//{'literal': 40, 'z': 8, 'op': 'literal'}
    instructions[576] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[577] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[578] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[579] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[580] = {5'd7, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'equal'}
    instructions[581] = {5'd6, 4'd0, 4'd8, 32'd585};//{'a': 8, 'label': 585, 'op': 'jmp_if_false'}
    instructions[582] = {5'd0, 4'd8, 4'd0, 32'd50};//{'literal': 50, 'z': 8, 'op': 'literal'}
    instructions[583] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[584] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[585] = {5'd6, 4'd0, 4'd8, 32'd588};//{'a': 8, 'label': 588, 'op': 'jmp_if_false'}
    instructions[586] = {5'd8, 4'd0, 4'd0, 32'd589};//{'label': 589, 'op': 'goto'}
    instructions[587] = {5'd8, 4'd0, 4'd0, 32'd588};//{'label': 588, 'op': 'goto'}
    instructions[588] = {5'd8, 4'd0, 4'd0, 32'd462};//{'label': 462, 'op': 'goto'}
    instructions[589] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[590] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[591] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[592] = {5'd1, 4'd8, 4'd4, 32'd2050};//{'a': 4, 'literal': 2050, 'z': 8, 'op': 'addl'}
    instructions[593] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[594] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[595] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[596] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[597] = {5'd7, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'equal'}
    instructions[598] = {5'd6, 4'd0, 4'd8, 32'd632};//{'a': 8, 'label': 632, 'op': 'jmp_if_false'}
    instructions[599] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[600] = {5'd0, 4'd2, 4'd0, 32'd1079};//{'literal': 1079, 'z': 2, 'op': 'literal'}
    instructions[601] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[602] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[603] = {5'd0, 4'd2, 4'd0, 32'd2704};//{'literal': 2704, 'z': 2, 'op': 'literal'}
    instructions[604] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[605] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[606] = {5'd0, 4'd2, 4'd0, 32'd2699};//{'literal': 2699, 'z': 2, 'op': 'literal'}
    instructions[607] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[608] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[609] = {5'd0, 4'd2, 4'd0, 32'd41};//{'literal': 41, 'z': 2, 'op': 'literal'}
    instructions[610] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[611] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[612] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[613] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[614] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[615] = {5'd1, 4'd8, 4'd4, 32'd1024};//{'a': 4, 'literal': 1024, 'z': 8, 'op': 'addl'}
    instructions[616] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[617] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[618] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[619] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[620] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[621] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[622] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[623] = {5'd3, 4'd6, 4'd0, 32'd4384};//{'z': 6, 'label': 4384, 'op': 'call'}
    instructions[624] = {5'd1, 4'd3, 4'd3, -32'd2};//{'a': 3, 'literal': -2, 'z': 3, 'op': 'addl'}
    instructions[625] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[626] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[627] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[628] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[629] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[630] = {5'd8, 4'd0, 4'd0, 32'd322};//{'label': 322, 'op': 'goto'}
    instructions[631] = {5'd8, 4'd0, 4'd0, 32'd632};//{'label': 632, 'op': 'goto'}
    instructions[632] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[633] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[634] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[635] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[636] = {5'd0, 4'd8, 4'd0, 32'd3};//{'literal': 3, 'z': 8, 'op': 'literal'}
    instructions[637] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[638] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[639] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[640] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[641] = {5'd3, 4'd6, 4'd0, 32'd1264};//{'z': 6, 'label': 1264, 'op': 'call'}
    instructions[642] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[643] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[644] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[645] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[646] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[647] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[648] = {5'd0, 4'd8, 4'd0, 32'd2723};//{'literal': 2723, 'z': 8, 'op': 'literal'}
    instructions[649] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[650] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[651] = {5'd0, 4'd2, 4'd0, 32'd2703};//{'literal': 2703, 'z': 2, 'op': 'literal'}
    instructions[652] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[653] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[654] = {5'd0, 4'd2, 4'd0, 32'd1079};//{'literal': 1079, 'z': 2, 'op': 'literal'}
    instructions[655] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[656] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[657] = {5'd0, 4'd2, 4'd0, 32'd2699};//{'literal': 2699, 'z': 2, 'op': 'literal'}
    instructions[658] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[659] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[660] = {5'd0, 4'd2, 4'd0, 32'd34};//{'literal': 34, 'z': 2, 'op': 'literal'}
    instructions[661] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[662] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[663] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[664] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[665] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[666] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[667] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[668] = {5'd3, 4'd6, 4'd0, 32'd5277};//{'z': 6, 'label': 5277, 'op': 'call'}
    instructions[669] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[670] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[671] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[672] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[673] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[674] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[675] = {5'd0, 4'd8, 4'd0, 32'd2703};//{'literal': 2703, 'z': 8, 'op': 'literal'}
    instructions[676] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[677] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[678] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[679] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[680] = {5'd0, 4'd8, 4'd0, 32'd2723};//{'literal': 2723, 'z': 8, 'op': 'literal'}
    instructions[681] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[682] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[683] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[684] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[685] = {5'd7, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'equal'}
    instructions[686] = {5'd6, 4'd0, 4'd8, 32'd741};//{'a': 8, 'label': 741, 'op': 'jmp_if_false'}
    instructions[687] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[688] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[689] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[690] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[691] = {5'd1, 4'd8, 4'd4, 32'd1024};//{'a': 4, 'literal': 1024, 'z': 8, 'op': 'addl'}
    instructions[692] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[693] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[694] = {5'd1, 4'd8, 4'd4, 32'd2048};//{'a': 4, 'literal': 2048, 'z': 8, 'op': 'addl'}
    instructions[695] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[696] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[697] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[698] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[699] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[700] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[701] = {5'd3, 4'd6, 4'd0, 32'd5467};//{'z': 6, 'label': 5467, 'op': 'call'}
    instructions[702] = {5'd1, 4'd3, 4'd3, -32'd2};//{'a': 3, 'literal': -2, 'z': 3, 'op': 'addl'}
    instructions[703] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[704] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[705] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[706] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[707] = {5'd0, 4'd2, 4'd0, 32'd2155};//{'literal': 2155, 'z': 2, 'op': 'literal'}
    instructions[708] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[709] = {5'd1, 4'd2, 4'd4, 32'd2049};//{'a': 4, 'literal': 2049, 'z': 2, 'op': 'addl'}
    instructions[710] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[711] = {5'd1, 4'd8, 4'd4, 32'd2049};//{'a': 4, 'literal': 2049, 'z': 8, 'op': 'addl'}
    instructions[712] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[713] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[714] = {5'd6, 4'd0, 4'd8, 32'd737};//{'a': 8, 'label': 737, 'op': 'jmp_if_false'}
    instructions[715] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[716] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[717] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[718] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[719] = {5'd1, 4'd8, 4'd4, 32'd1024};//{'a': 4, 'literal': 1024, 'z': 8, 'op': 'addl'}
    instructions[720] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[721] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[722] = {5'd1, 4'd8, 4'd4, 32'd2049};//{'a': 4, 'literal': 2049, 'z': 8, 'op': 'addl'}
    instructions[723] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[724] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[725] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[726] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[727] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[728] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[729] = {5'd3, 4'd6, 4'd0, 32'd4384};//{'z': 6, 'label': 4384, 'op': 'call'}
    instructions[730] = {5'd1, 4'd3, 4'd3, -32'd2};//{'a': 3, 'literal': -2, 'z': 3, 'op': 'addl'}
    instructions[731] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[732] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[733] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[734] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[735] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[736] = {5'd8, 4'd0, 4'd0, 32'd737};//{'label': 737, 'op': 'goto'}
    instructions[737] = {5'd0, 4'd8, 4'd0, 32'd10000};//{'literal': 10000, 'z': 8, 'op': 'literal'}
    instructions[738] = {5'd1, 4'd2, 4'd4, 32'd2053};//{'a': 4, 'literal': 2053, 'z': 2, 'op': 'addl'}
    instructions[739] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[740] = {5'd8, 4'd0, 4'd0, 32'd815};//{'label': 815, 'op': 'goto'}
    instructions[741] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[742] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[743] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[744] = {5'd1, 4'd8, 4'd4, 32'd2053};//{'a': 4, 'literal': 2053, 'z': 8, 'op': 'addl'}
    instructions[745] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[746] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[747] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[748] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[749] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[750] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[751] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[752] = {5'd1, 4'd8, 4'd4, 32'd2053};//{'a': 4, 'literal': 2053, 'z': 8, 'op': 'addl'}
    instructions[753] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[754] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[755] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[756] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[757] = {5'd10, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'subtract'}
    instructions[758] = {5'd1, 4'd2, 4'd4, 32'd2053};//{'a': 4, 'literal': 2053, 'z': 2, 'op': 'addl'}
    instructions[759] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[760] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[761] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[762] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[763] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[764] = {5'd7, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'equal'}
    instructions[765] = {5'd6, 4'd0, 4'd8, 32'd815};//{'a': 8, 'label': 815, 'op': 'jmp_if_false'}
    instructions[766] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[767] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[768] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[769] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[770] = {5'd1, 4'd8, 4'd4, 32'd1024};//{'a': 4, 'literal': 1024, 'z': 8, 'op': 'addl'}
    instructions[771] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[772] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[773] = {5'd1, 4'd8, 4'd4, 32'd2048};//{'a': 4, 'literal': 2048, 'z': 8, 'op': 'addl'}
    instructions[774] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[775] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[776] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[777] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[778] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[779] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[780] = {5'd3, 4'd6, 4'd0, 32'd5467};//{'z': 6, 'label': 5467, 'op': 'call'}
    instructions[781] = {5'd1, 4'd3, 4'd3, -32'd2};//{'a': 3, 'literal': -2, 'z': 3, 'op': 'addl'}
    instructions[782] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[783] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[784] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[785] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[786] = {5'd0, 4'd2, 4'd0, 32'd2155};//{'literal': 2155, 'z': 2, 'op': 'literal'}
    instructions[787] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[788] = {5'd1, 4'd2, 4'd4, 32'd2049};//{'a': 4, 'literal': 2049, 'z': 2, 'op': 'addl'}
    instructions[789] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[790] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[791] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[792] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[793] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[794] = {5'd1, 4'd8, 4'd4, 32'd1024};//{'a': 4, 'literal': 1024, 'z': 8, 'op': 'addl'}
    instructions[795] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[796] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[797] = {5'd1, 4'd8, 4'd4, 32'd2049};//{'a': 4, 'literal': 2049, 'z': 8, 'op': 'addl'}
    instructions[798] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[799] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[800] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[801] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[802] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[803] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[804] = {5'd3, 4'd6, 4'd0, 32'd4384};//{'z': 6, 'label': 4384, 'op': 'call'}
    instructions[805] = {5'd1, 4'd3, 4'd3, -32'd2};//{'a': 3, 'literal': -2, 'z': 3, 'op': 'addl'}
    instructions[806] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[807] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[808] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[809] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[810] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[811] = {5'd0, 4'd8, 4'd0, 32'd10000};//{'literal': 10000, 'z': 8, 'op': 'literal'}
    instructions[812] = {5'd1, 4'd2, 4'd4, 32'd2053};//{'a': 4, 'literal': 2053, 'z': 2, 'op': 'addl'}
    instructions[813] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[814] = {5'd8, 4'd0, 4'd0, 32'd815};//{'label': 815, 'op': 'goto'}
    instructions[815] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[816] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[817] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[818] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[819] = {5'd1, 4'd8, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 8, 'op': 'addl'}
    instructions[820] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[821] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[822] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[823] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[824] = {5'd3, 4'd6, 4'd0, 32'd1352};//{'z': 6, 'label': 1352, 'op': 'call'}
    instructions[825] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[826] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[827] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[828] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[829] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[830] = {5'd0, 4'd2, 4'd0, 32'd2701};//{'literal': 2701, 'z': 2, 'op': 'literal'}
    instructions[831] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[832] = {5'd6, 4'd0, 4'd8, 32'd842};//{'a': 8, 'label': 842, 'op': 'jmp_if_false'}
    instructions[833] = {5'd0, 4'd8, 4'd0, 32'd80};//{'literal': 80, 'z': 8, 'op': 'literal'}
    instructions[834] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[835] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[836] = {5'd0, 4'd8, 4'd0, 32'd2726};//{'literal': 2726, 'z': 8, 'op': 'literal'}
    instructions[837] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[838] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[839] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[840] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[841] = {5'd7, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'equal'}
    instructions[842] = {5'd6, 4'd0, 4'd8, 32'd854};//{'a': 8, 'label': 854, 'op': 'jmp_if_false'}
    instructions[843] = {5'd0, 4'd8, 4'd0, 32'd1078};//{'literal': 1078, 'z': 8, 'op': 'literal'}
    instructions[844] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[845] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[846] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[847] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[848] = {5'd0, 4'd8, 4'd0, 32'd40};//{'literal': 40, 'z': 8, 'op': 'literal'}
    instructions[849] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[850] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[851] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[852] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[853] = {5'd7, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'equal'}
    instructions[854] = {5'd6, 4'd0, 4'd8, 32'd972};//{'a': 8, 'label': 972, 'op': 'jmp_if_false'}
    instructions[855] = {5'd0, 4'd8, 4'd0, 32'd46};//{'literal': 46, 'z': 8, 'op': 'literal'}
    instructions[856] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[857] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[858] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[859] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[860] = {5'd0, 4'd8, 4'd0, 32'd2};//{'literal': 2, 'z': 8, 'op': 'literal'}
    instructions[861] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[862] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[863] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[864] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[865] = {5'd7, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'equal'}
    instructions[866] = {5'd6, 4'd0, 4'd8, 32'd929};//{'a': 8, 'label': 929, 'op': 'jmp_if_false'}
    instructions[867] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[868] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[869] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[870] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[871] = {5'd1, 4'd8, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 8, 'op': 'addl'}
    instructions[872] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[873] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[874] = {5'd0, 4'd8, 4'd0, 32'd48};//{'literal': 48, 'z': 8, 'op': 'literal'}
    instructions[875] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[876] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[877] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[878] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[879] = {5'd0, 4'd8, 4'd0, 32'd1122};//{'literal': 1122, 'z': 8, 'op': 'literal'}
    instructions[880] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[881] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[882] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[883] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[884] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[885] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[886] = {5'd3, 4'd6, 4'd0, 32'd5721};//{'z': 6, 'label': 5721, 'op': 'call'}
    instructions[887] = {5'd1, 4'd3, 4'd3, -32'd3};//{'a': 3, 'literal': -3, 'z': 3, 'op': 'addl'}
    instructions[888] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[889] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[890] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[891] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[892] = {5'd0, 4'd2, 4'd0, 32'd2700};//{'literal': 2700, 'z': 2, 'op': 'literal'}
    instructions[893] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[894] = {5'd6, 4'd0, 4'd8, 32'd928};//{'a': 8, 'label': 928, 'op': 'jmp_if_false'}
    instructions[895] = {5'd0, 4'd8, 4'd0, 32'd1122};//{'literal': 1122, 'z': 8, 'op': 'literal'}
    instructions[896] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[897] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[898] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[899] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[900] = {5'd0, 4'd8, 4'd0, 32'd2};//{'literal': 2, 'z': 8, 'op': 'literal'}
    instructions[901] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[902] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[903] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[904] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[905] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[906] = {5'd0, 4'd2, 4'd0, 32'd46};//{'literal': 46, 'z': 2, 'op': 'literal'}
    instructions[907] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[908] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[909] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[910] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[911] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[912] = {5'd1, 4'd8, 4'd4, 32'd1024};//{'a': 4, 'literal': 1024, 'z': 8, 'op': 'addl'}
    instructions[913] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[914] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[915] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[916] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[917] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[918] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[919] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[920] = {5'd3, 4'd6, 4'd0, 32'd4384};//{'z': 6, 'label': 4384, 'op': 'call'}
    instructions[921] = {5'd1, 4'd3, 4'd3, -32'd2};//{'a': 3, 'literal': -2, 'z': 3, 'op': 'addl'}
    instructions[922] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[923] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[924] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[925] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[926] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[927] = {5'd8, 4'd0, 4'd0, 32'd928};//{'label': 928, 'op': 'goto'}
    instructions[928] = {5'd8, 4'd0, 4'd0, 32'd929};//{'label': 929, 'op': 'goto'}
    instructions[929] = {5'd0, 4'd8, 4'd0, 32'd50};//{'literal': 50, 'z': 8, 'op': 'literal'}
    instructions[930] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[931] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[932] = {5'd6, 4'd0, 4'd8, 32'd965};//{'a': 8, 'label': 965, 'op': 'jmp_if_false'}
    instructions[933] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[934] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[935] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[936] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[937] = {5'd0, 4'd8, 4'd0, 32'd2703};//{'literal': 2703, 'z': 8, 'op': 'literal'}
    instructions[938] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[939] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[940] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[941] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[942] = {5'd0, 4'd8, 4'd0, 32'd2723};//{'literal': 2723, 'z': 8, 'op': 'literal'}
    instructions[943] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[944] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[945] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[946] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[947] = {5'd10, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'subtract'}
    instructions[948] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[949] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[950] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[951] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[952] = {5'd3, 4'd6, 4'd0, 32'd5945};//{'z': 6, 'label': 5945, 'op': 'call'}
    instructions[953] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[954] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[955] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[956] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[957] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[958] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[959] = {5'd0, 4'd8, 4'd0, 32'd2723};//{'literal': 2723, 'z': 8, 'op': 'literal'}
    instructions[960] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[961] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[962] = {5'd0, 4'd2, 4'd0, 32'd2703};//{'literal': 2703, 'z': 2, 'op': 'literal'}
    instructions[963] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[964] = {5'd8, 4'd0, 4'd0, 32'd965};//{'label': 965, 'op': 'goto'}
    instructions[965] = {5'd0, 4'd8, 4'd0, 32'd2722};//{'literal': 2722, 'z': 8, 'op': 'literal'}
    instructions[966] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[967] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[968] = {5'd6, 4'd0, 4'd8, 32'd971};//{'a': 8, 'label': 971, 'op': 'jmp_if_false'}
    instructions[969] = {5'd8, 4'd0, 4'd0, 32'd973};//{'label': 973, 'op': 'goto'}
    instructions[970] = {5'd8, 4'd0, 4'd0, 32'd971};//{'label': 971, 'op': 'goto'}
    instructions[971] = {5'd8, 4'd0, 4'd0, 32'd972};//{'label': 972, 'op': 'goto'}
    instructions[972] = {5'd8, 4'd0, 4'd0, 32'd662};//{'label': 662, 'op': 'goto'}
    instructions[973] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[974] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[975] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[976] = {5'd1, 4'd8, 4'd4, 32'd2050};//{'a': 4, 'literal': 2050, 'z': 8, 'op': 'addl'}
    instructions[977] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[978] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[979] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[980] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[981] = {5'd7, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'equal'}
    instructions[982] = {5'd6, 4'd0, 4'd8, 32'd1019};//{'a': 8, 'label': 1019, 'op': 'jmp_if_false'}
    instructions[983] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[984] = {5'd0, 4'd2, 4'd0, 32'd34};//{'literal': 34, 'z': 2, 'op': 'literal'}
    instructions[985] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[986] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[987] = {5'd0, 4'd2, 4'd0, 32'd1079};//{'literal': 1079, 'z': 2, 'op': 'literal'}
    instructions[988] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[989] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[990] = {5'd0, 4'd2, 4'd0, 32'd2704};//{'literal': 2704, 'z': 2, 'op': 'literal'}
    instructions[991] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[992] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[993] = {5'd0, 4'd2, 4'd0, 32'd2699};//{'literal': 2699, 'z': 2, 'op': 'literal'}
    instructions[994] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[995] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[996] = {5'd0, 4'd2, 4'd0, 32'd41};//{'literal': 41, 'z': 2, 'op': 'literal'}
    instructions[997] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[998] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[999] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1000] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[1001] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1002] = {5'd1, 4'd8, 4'd4, 32'd1024};//{'a': 4, 'literal': 1024, 'z': 8, 'op': 'addl'}
    instructions[1003] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1004] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1005] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[1006] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1007] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1008] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[1009] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[1010] = {5'd3, 4'd6, 4'd0, 32'd4384};//{'z': 6, 'label': 4384, 'op': 'call'}
    instructions[1011] = {5'd1, 4'd3, 4'd3, -32'd2};//{'a': 3, 'literal': -2, 'z': 3, 'op': 'addl'}
    instructions[1012] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1013] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[1014] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1015] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[1016] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[1017] = {5'd8, 4'd0, 4'd0, 32'd322};//{'label': 322, 'op': 'goto'}
    instructions[1018] = {5'd8, 4'd0, 4'd0, 32'd1019};//{'label': 1019, 'op': 'goto'}
    instructions[1019] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[1020] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1021] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[1022] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1023] = {5'd0, 4'd8, 4'd0, 32'd1110};//{'literal': 1110, 'z': 8, 'op': 'literal'}
    instructions[1024] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1025] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1026] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[1027] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[1028] = {5'd3, 4'd6, 4'd0, 32'd1264};//{'z': 6, 'label': 1264, 'op': 'call'}
    instructions[1029] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1030] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1031] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[1032] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1033] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[1034] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[1035] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[1036] = {5'd0, 4'd2, 4'd0, 32'd34};//{'literal': 34, 'z': 2, 'op': 'literal'}
    instructions[1037] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1038] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[1039] = {5'd0, 4'd2, 4'd0, 32'd2704};//{'literal': 2704, 'z': 2, 'op': 'literal'}
    instructions[1040] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1041] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[1042] = {5'd0, 4'd2, 4'd0, 32'd2699};//{'literal': 2699, 'z': 2, 'op': 'literal'}
    instructions[1043] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1044] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[1045] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1046] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1047] = {5'd0, 4'd8, 4'd0, 32'd2};//{'literal': 2, 'z': 8, 'op': 'literal'}
    instructions[1048] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1049] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1050] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1051] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1052] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[1053] = {5'd0, 4'd2, 4'd0, 32'd46};//{'literal': 46, 'z': 2, 'op': 'literal'}
    instructions[1054] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1055] = {5'd0, 4'd8, 4'd0, 32'd10000};//{'literal': 10000, 'z': 8, 'op': 'literal'}
    instructions[1056] = {5'd1, 4'd2, 4'd4, 32'd2050};//{'a': 4, 'literal': 2050, 'z': 2, 'op': 'addl'}
    instructions[1057] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1058] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[1059] = {5'd1, 4'd2, 4'd4, 32'd2052};//{'a': 4, 'literal': 2052, 'z': 2, 'op': 'addl'}
    instructions[1060] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1061] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[1062] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1063] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1064] = {5'd1, 4'd8, 4'd4, 32'd2052};//{'a': 4, 'literal': 2052, 'z': 8, 'op': 'addl'}
    instructions[1065] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1066] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1067] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1068] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1069] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[1070] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1071] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1072] = {5'd1, 4'd8, 4'd4, 32'd2052};//{'a': 4, 'literal': 2052, 'z': 8, 'op': 'addl'}
    instructions[1073] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1074] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1075] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1076] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1077] = {5'd10, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'subtract'}
    instructions[1078] = {5'd1, 4'd2, 4'd4, 32'd2052};//{'a': 4, 'literal': 2052, 'z': 2, 'op': 'addl'}
    instructions[1079] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1080] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1081] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[1082] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1083] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1084] = {5'd7, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'equal'}
    instructions[1085] = {5'd6, 4'd0, 4'd8, 32'd1136};//{'a': 8, 'label': 1136, 'op': 'jmp_if_false'}
    instructions[1086] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[1087] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1088] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[1089] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1090] = {5'd1, 4'd8, 4'd4, 32'd1024};//{'a': 4, 'literal': 1024, 'z': 8, 'op': 'addl'}
    instructions[1091] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1092] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1093] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[1094] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1095] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1096] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[1097] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[1098] = {5'd3, 4'd6, 4'd0, 32'd4384};//{'z': 6, 'label': 4384, 'op': 'call'}
    instructions[1099] = {5'd1, 4'd3, 4'd3, -32'd2};//{'a': 3, 'literal': -2, 'z': 3, 'op': 'addl'}
    instructions[1100] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1101] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[1102] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1103] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[1104] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[1105] = {5'd0, 4'd8, 4'd0, 32'd10};//{'literal': 10, 'z': 8, 'op': 'literal'}
    instructions[1106] = {5'd1, 4'd2, 4'd4, 32'd2052};//{'a': 4, 'literal': 2052, 'z': 2, 'op': 'addl'}
    instructions[1107] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1108] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[1109] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1110] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1111] = {5'd1, 4'd8, 4'd4, 32'd2050};//{'a': 4, 'literal': 2050, 'z': 8, 'op': 'addl'}
    instructions[1112] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1113] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1114] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1115] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1116] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[1117] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1118] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1119] = {5'd1, 4'd8, 4'd4, 32'd2050};//{'a': 4, 'literal': 2050, 'z': 8, 'op': 'addl'}
    instructions[1120] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1121] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1122] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1123] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1124] = {5'd10, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'subtract'}
    instructions[1125] = {5'd1, 4'd2, 4'd4, 32'd2050};//{'a': 4, 'literal': 2050, 'z': 2, 'op': 'addl'}
    instructions[1126] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1127] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1128] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[1129] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1130] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1131] = {5'd7, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'equal'}
    instructions[1132] = {5'd6, 4'd0, 4'd8, 32'd1135};//{'a': 8, 'label': 1135, 'op': 'jmp_if_false'}
    instructions[1133] = {5'd8, 4'd0, 4'd0, 32'd1217};//{'label': 1217, 'op': 'goto'}
    instructions[1134] = {5'd8, 4'd0, 4'd0, 32'd1135};//{'label': 1135, 'op': 'goto'}
    instructions[1135] = {5'd8, 4'd0, 4'd0, 32'd1136};//{'label': 1136, 'op': 'goto'}
    instructions[1136] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[1137] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1138] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[1139] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1140] = {5'd1, 4'd8, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 8, 'op': 'addl'}
    instructions[1141] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1142] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1143] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[1144] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[1145] = {5'd3, 4'd6, 4'd0, 32'd1352};//{'z': 6, 'label': 1352, 'op': 'call'}
    instructions[1146] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1147] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1148] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[1149] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1150] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[1151] = {5'd0, 4'd2, 4'd0, 32'd2701};//{'literal': 2701, 'z': 2, 'op': 'literal'}
    instructions[1152] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1153] = {5'd1, 4'd2, 4'd4, 32'd2051};//{'a': 4, 'literal': 2051, 'z': 2, 'op': 'addl'}
    instructions[1154] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1155] = {5'd1, 4'd8, 4'd4, 32'd2051};//{'a': 4, 'literal': 2051, 'z': 8, 'op': 'addl'}
    instructions[1156] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1157] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1158] = {5'd6, 4'd0, 4'd8, 32'd1168};//{'a': 8, 'label': 1168, 'op': 'jmp_if_false'}
    instructions[1159] = {5'd0, 4'd8, 4'd0, 32'd80};//{'literal': 80, 'z': 8, 'op': 'literal'}
    instructions[1160] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1161] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1162] = {5'd0, 4'd8, 4'd0, 32'd2726};//{'literal': 2726, 'z': 8, 'op': 'literal'}
    instructions[1163] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1164] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1165] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1166] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1167] = {5'd7, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'equal'}
    instructions[1168] = {5'd6, 4'd0, 4'd8, 32'd1180};//{'a': 8, 'label': 1180, 'op': 'jmp_if_false'}
    instructions[1169] = {5'd0, 4'd8, 4'd0, 32'd1078};//{'literal': 1078, 'z': 8, 'op': 'literal'}
    instructions[1170] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1171] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1172] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1173] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1174] = {5'd0, 4'd8, 4'd0, 32'd40};//{'literal': 40, 'z': 8, 'op': 'literal'}
    instructions[1175] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1176] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1177] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1178] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1179] = {5'd7, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'equal'}
    instructions[1180] = {5'd6, 4'd0, 4'd8, 32'd1184};//{'a': 8, 'label': 1184, 'op': 'jmp_if_false'}
    instructions[1181] = {5'd0, 4'd8, 4'd0, 32'd50};//{'literal': 50, 'z': 8, 'op': 'literal'}
    instructions[1182] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1183] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1184] = {5'd6, 4'd0, 4'd8, 32'd1187};//{'a': 8, 'label': 1187, 'op': 'jmp_if_false'}
    instructions[1185] = {5'd8, 4'd0, 4'd0, 32'd1217};//{'label': 1217, 'op': 'goto'}
    instructions[1186] = {5'd8, 4'd0, 4'd0, 32'd1187};//{'label': 1187, 'op': 'goto'}
    instructions[1187] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[1188] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1189] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1190] = {5'd1, 4'd8, 4'd4, 32'd2050};//{'a': 4, 'literal': 2050, 'z': 8, 'op': 'addl'}
    instructions[1191] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1192] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1193] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1194] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1195] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[1196] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1197] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1198] = {5'd1, 4'd8, 4'd4, 32'd2050};//{'a': 4, 'literal': 2050, 'z': 8, 'op': 'addl'}
    instructions[1199] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1200] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1201] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1202] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1203] = {5'd10, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'subtract'}
    instructions[1204] = {5'd1, 4'd2, 4'd4, 32'd2050};//{'a': 4, 'literal': 2050, 'z': 2, 'op': 'addl'}
    instructions[1205] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1206] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1207] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[1208] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1209] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1210] = {5'd7, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'equal'}
    instructions[1211] = {5'd6, 4'd0, 4'd8, 32'd1214};//{'a': 8, 'label': 1214, 'op': 'jmp_if_false'}
    instructions[1212] = {5'd8, 4'd0, 4'd0, 32'd1217};//{'label': 1217, 'op': 'goto'}
    instructions[1213] = {5'd8, 4'd0, 4'd0, 32'd1214};//{'label': 1214, 'op': 'goto'}
    instructions[1214] = {5'd0, 4'd8, 4'd0, 32'd5000};//{'literal': 5000, 'z': 8, 'op': 'literal'}
    instructions[1215] = {5'd11, 4'd0, 4'd8, 32'd0};//{'a': 8, 'op': 'wait_clocks'}
    instructions[1216] = {5'd8, 4'd0, 4'd0, 32'd1061};//{'label': 1061, 'op': 'goto'}
    instructions[1217] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[1218] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1219] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1220] = {5'd1, 4'd8, 4'd4, 32'd2050};//{'a': 4, 'literal': 2050, 'z': 8, 'op': 'addl'}
    instructions[1221] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1222] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1223] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1224] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1225] = {5'd7, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'equal'}
    instructions[1226] = {5'd6, 4'd0, 4'd8, 32'd1260};//{'a': 8, 'label': 1260, 'op': 'jmp_if_false'}
    instructions[1227] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[1228] = {5'd0, 4'd2, 4'd0, 32'd1079};//{'literal': 1079, 'z': 2, 'op': 'literal'}
    instructions[1229] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1230] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[1231] = {5'd0, 4'd2, 4'd0, 32'd2704};//{'literal': 2704, 'z': 2, 'op': 'literal'}
    instructions[1232] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1233] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[1234] = {5'd0, 4'd2, 4'd0, 32'd2699};//{'literal': 2699, 'z': 2, 'op': 'literal'}
    instructions[1235] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1236] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[1237] = {5'd0, 4'd2, 4'd0, 32'd41};//{'literal': 41, 'z': 2, 'op': 'literal'}
    instructions[1238] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1239] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[1240] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1241] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[1242] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1243] = {5'd1, 4'd8, 4'd4, 32'd1024};//{'a': 4, 'literal': 1024, 'z': 8, 'op': 'addl'}
    instructions[1244] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1245] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1246] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[1247] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1248] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1249] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[1250] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[1251] = {5'd3, 4'd6, 4'd0, 32'd4384};//{'z': 6, 'label': 4384, 'op': 'call'}
    instructions[1252] = {5'd1, 4'd3, 4'd3, -32'd2};//{'a': 3, 'literal': -2, 'z': 3, 'op': 'addl'}
    instructions[1253] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1254] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[1255] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1256] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[1257] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[1258] = {5'd8, 4'd0, 4'd0, 32'd322};//{'label': 322, 'op': 'goto'}
    instructions[1259] = {5'd8, 4'd0, 4'd0, 32'd1260};//{'label': 1260, 'op': 'goto'}
    instructions[1260] = {5'd8, 4'd0, 4'd0, 32'd322};//{'label': 322, 'op': 'goto'}
    instructions[1261] = {5'd1, 4'd3, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[1262] = {5'd1, 4'd4, 4'd7, 32'd0};//{'a': 7, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[1263] = {5'd12, 4'd0, 4'd6, 32'd0};//{'a': 6, 'op': 'return'}
    instructions[1264] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[1265] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[1266] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1267] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[1268] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1269] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[1270] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[1271] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1272] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1273] = {5'd0, 4'd8, 4'd0, 32'd47};//{'literal': 47, 'z': 8, 'op': 'literal'}
    instructions[1274] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1275] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1276] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1277] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1278] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[1279] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[1280] = {5'd3, 4'd6, 4'd0, 32'd1290};//{'z': 6, 'label': 1290, 'op': 'call'}
    instructions[1281] = {5'd1, 4'd3, 4'd3, -32'd2};//{'a': 3, 'literal': -2, 'z': 3, 'op': 'addl'}
    instructions[1282] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1283] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[1284] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1285] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[1286] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[1287] = {5'd1, 4'd3, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[1288] = {5'd1, 4'd4, 4'd7, 32'd0};//{'a': 7, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[1289] = {5'd12, 4'd0, 4'd6, 32'd0};//{'a': 6, 'op': 'return'}
    instructions[1290] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1291] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[1292] = {5'd1, 4'd2, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1293] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1294] = {5'd1, 4'd8, 4'd4, -32'd2};//{'a': 4, 'literal': -2, 'z': 8, 'op': 'addl'}
    instructions[1295] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[1296] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1297] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1298] = {5'd1, 4'd8, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 8, 'op': 'addl'}
    instructions[1299] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1300] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1301] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1302] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[1303] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[1304] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1305] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1306] = {5'd6, 4'd0, 4'd8, 32'd1347};//{'a': 8, 'label': 1347, 'op': 'jmp_if_false'}
    instructions[1307] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[1308] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1309] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1310] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1311] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1312] = {5'd1, 4'd8, 4'd4, -32'd2};//{'a': 4, 'literal': -2, 'z': 8, 'op': 'addl'}
    instructions[1313] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[1314] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1315] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1316] = {5'd1, 4'd8, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 8, 'op': 'addl'}
    instructions[1317] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1318] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1319] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1320] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[1321] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[1322] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1323] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1324] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1325] = {5'd5, 4'd0, 4'd3, 32'd0};//{'a': 3, 'z': 0, 'op': 'load'}
    instructions[1326] = {5'd13, 4'd0, 4'd0, 32'd8};//{'a': 0, 'b': 8, 'op': 'write'}
    instructions[1327] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[1328] = {5'd1, 4'd8, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 8, 'op': 'addl'}
    instructions[1329] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1330] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1331] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1332] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1333] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[1334] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1335] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1336] = {5'd1, 4'd8, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 8, 'op': 'addl'}
    instructions[1337] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1338] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1339] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1340] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1341] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[1342] = {5'd1, 4'd2, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1343] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1344] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1345] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[1346] = {5'd8, 4'd0, 4'd0, 32'd1348};//{'label': 1348, 'op': 'goto'}
    instructions[1347] = {5'd8, 4'd0, 4'd0, 32'd1349};//{'label': 1349, 'op': 'goto'}
    instructions[1348] = {5'd8, 4'd0, 4'd0, 32'd1294};//{'label': 1294, 'op': 'goto'}
    instructions[1349] = {5'd1, 4'd3, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[1350] = {5'd1, 4'd4, 4'd7, 32'd0};//{'a': 7, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[1351] = {5'd12, 4'd0, 4'd6, 32'd0};//{'a': 6, 'op': 'return'}
    instructions[1352] = {5'd1, 4'd3, 4'd3, 32'd7};//{'a': 3, 'literal': 7, 'z': 3, 'op': 'addl'}
    instructions[1353] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[1354] = {5'd1, 4'd2, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1355] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1356] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[1357] = {5'd1, 4'd2, 4'd4, 32'd1};//{'a': 4, 'literal': 1, 'z': 2, 'op': 'addl'}
    instructions[1358] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1359] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[1360] = {5'd1, 4'd2, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 2, 'op': 'addl'}
    instructions[1361] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1362] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[1363] = {5'd1, 4'd2, 4'd4, 32'd3};//{'a': 4, 'literal': 3, 'z': 2, 'op': 'addl'}
    instructions[1364] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1365] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[1366] = {5'd1, 4'd2, 4'd4, 32'd4};//{'a': 4, 'literal': 4, 'z': 2, 'op': 'addl'}
    instructions[1367] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1368] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[1369] = {5'd1, 4'd2, 4'd4, 32'd5};//{'a': 4, 'literal': 5, 'z': 2, 'op': 'addl'}
    instructions[1370] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1371] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[1372] = {5'd1, 4'd2, 4'd4, 32'd6};//{'a': 4, 'literal': 6, 'z': 2, 'op': 'addl'}
    instructions[1373] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1374] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[1375] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1376] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[1377] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1378] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[1379] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[1380] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1381] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1382] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[1383] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[1384] = {5'd3, 4'd6, 4'd0, 32'd1862};//{'z': 6, 'label': 1862, 'op': 'call'}
    instructions[1385] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1386] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1387] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[1388] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1389] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[1390] = {5'd0, 4'd2, 4'd0, 32'd42};//{'literal': 42, 'z': 2, 'op': 'literal'}
    instructions[1391] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1392] = {5'd1, 4'd2, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1393] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1394] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[1395] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1396] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1397] = {5'd0, 4'd8, 4'd0, 32'd15};//{'literal': 15, 'z': 8, 'op': 'literal'}
    instructions[1398] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1399] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1400] = {5'd0, 4'd8, 4'd0, 32'd8};//{'literal': 8, 'z': 8, 'op': 'literal'}
    instructions[1401] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1402] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1403] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[1404] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[1405] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1406] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1407] = {5'd0, 4'd8, 4'd0, 32'd7};//{'literal': 7, 'z': 8, 'op': 'literal'}
    instructions[1408] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1409] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[1410] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[1411] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1412] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1413] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1414] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1415] = {5'd14, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'unsigned_shift_right'}
    instructions[1416] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1417] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1418] = {5'd15, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'and'}
    instructions[1419] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1420] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1421] = {5'd16, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'shift_left'}
    instructions[1422] = {5'd1, 4'd2, 4'd4, 32'd1};//{'a': 4, 'literal': 1, 'z': 2, 'op': 'addl'}
    instructions[1423] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1424] = {5'd0, 4'd8, 4'd0, 32'd7};//{'literal': 7, 'z': 8, 'op': 'literal'}
    instructions[1425] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1426] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1427] = {5'd1, 4'd8, 4'd4, 32'd1};//{'a': 4, 'literal': 1, 'z': 8, 'op': 'addl'}
    instructions[1428] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1429] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1430] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1431] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1432] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[1433] = {5'd1, 4'd2, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 2, 'op': 'addl'}
    instructions[1434] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1435] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[1436] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[1437] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1438] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1439] = {5'd0, 4'd8, 4'd0, 32'd8};//{'literal': 8, 'z': 8, 'op': 'literal'}
    instructions[1440] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1441] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[1442] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[1443] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1444] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1445] = {5'd1, 4'd2, 4'd4, 32'd3};//{'a': 4, 'literal': 3, 'z': 2, 'op': 'addl'}
    instructions[1446] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1447] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[1448] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1449] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1450] = {5'd1, 4'd8, 4'd4, 32'd1};//{'a': 4, 'literal': 1, 'z': 8, 'op': 'addl'}
    instructions[1451] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1452] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1453] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1454] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1455] = {5'd16, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'shift_left'}
    instructions[1456] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1457] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1458] = {5'd1, 4'd8, 4'd4, 32'd3};//{'a': 4, 'literal': 3, 'z': 8, 'op': 'addl'}
    instructions[1459] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1460] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1461] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1462] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1463] = {5'd10, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'subtract'}
    instructions[1464] = {5'd1, 4'd2, 4'd4, 32'd4};//{'a': 4, 'literal': 4, 'z': 2, 'op': 'addl'}
    instructions[1465] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1466] = {5'd0, 4'd8, 4'd0, 32'd10};//{'literal': 10, 'z': 8, 'op': 'literal'}
    instructions[1467] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1468] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1469] = {5'd0, 4'd8, 4'd0, 32'd61440};//{'literal': 61440, 'z': 8, 'op': 'literal'}
    instructions[1470] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1471] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1472] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[1473] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[1474] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1475] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1476] = {5'd0, 4'd8, 4'd0, 32'd6};//{'literal': 6, 'z': 8, 'op': 'literal'}
    instructions[1477] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1478] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1479] = {5'd1, 4'd8, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 8, 'op': 'addl'}
    instructions[1480] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1481] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1482] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1483] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1484] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[1485] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1486] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[1487] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[1488] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1489] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1490] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1491] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1492] = {5'd15, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'and'}
    instructions[1493] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1494] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1495] = {5'd14, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'unsigned_shift_right'}
    instructions[1496] = {5'd1, 4'd2, 4'd4, 32'd6};//{'a': 4, 'literal': 6, 'z': 2, 'op': 'addl'}
    instructions[1497] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1498] = {5'd1, 4'd8, 4'd4, 32'd6};//{'a': 4, 'literal': 6, 'z': 8, 'op': 'addl'}
    instructions[1499] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1500] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1501] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1502] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1503] = {5'd1, 4'd8, 4'd4, 32'd4};//{'a': 4, 'literal': 4, 'z': 8, 'op': 'addl'}
    instructions[1504] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1505] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1506] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1507] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1508] = {5'd10, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'subtract'}
    instructions[1509] = {5'd0, 4'd2, 4'd0, 32'd1122};//{'literal': 1122, 'z': 2, 'op': 'literal'}
    instructions[1510] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1511] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[1512] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1513] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1514] = {5'd1, 4'd8, 4'd4, 32'd6};//{'a': 4, 'literal': 6, 'z': 8, 'op': 'addl'}
    instructions[1515] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1516] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1517] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1518] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1519] = {5'd14, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'unsigned_shift_right'}
    instructions[1520] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1521] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1522] = {5'd1, 4'd8, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 8, 'op': 'addl'}
    instructions[1523] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1524] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1525] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1526] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1527] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[1528] = {5'd0, 4'd2, 4'd0, 32'd48};//{'literal': 48, 'z': 2, 'op': 'literal'}
    instructions[1529] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1530] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[1531] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[1532] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1533] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1534] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[1535] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1536] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1537] = {5'd1, 4'd8, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 8, 'op': 'addl'}
    instructions[1538] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1539] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1540] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1541] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1542] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[1543] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1544] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[1545] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[1546] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1547] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1548] = {5'd0, 4'd2, 4'd0, 32'd40};//{'literal': 40, 'z': 2, 'op': 'literal'}
    instructions[1549] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1550] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[1551] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[1552] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1553] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1554] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[1555] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1556] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1557] = {5'd1, 4'd8, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 8, 'op': 'addl'}
    instructions[1558] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1559] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1560] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1561] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1562] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[1563] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1564] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[1565] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[1566] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1567] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1568] = {5'd0, 4'd2, 4'd0, 32'd2726};//{'literal': 2726, 'z': 2, 'op': 'literal'}
    instructions[1569] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1570] = {5'd0, 4'd8, 4'd0, 32'd16};//{'literal': 16, 'z': 8, 'op': 'literal'}
    instructions[1571] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1572] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1573] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[1574] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[1575] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1576] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1577] = {5'd0, 4'd8, 4'd0, 32'd2};//{'literal': 2, 'z': 8, 'op': 'literal'}
    instructions[1578] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1579] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1580] = {5'd1, 4'd8, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 8, 'op': 'addl'}
    instructions[1581] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1582] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1583] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1584] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1585] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[1586] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1587] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[1588] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[1589] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1590] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1591] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1592] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1593] = {5'd16, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'shift_left'}
    instructions[1594] = {5'd0, 4'd2, 4'd0, 32'd2};//{'literal': 2, 'z': 2, 'op': 'literal'}
    instructions[1595] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1596] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[1597] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[1598] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1599] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1600] = {5'd0, 4'd8, 4'd0, 32'd3};//{'literal': 3, 'z': 8, 'op': 'literal'}
    instructions[1601] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1602] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1603] = {5'd1, 4'd8, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 8, 'op': 'addl'}
    instructions[1604] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1605] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1606] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1607] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1608] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[1609] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1610] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[1611] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[1612] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1613] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1614] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1615] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1616] = {5'd0, 4'd8, 4'd0, 32'd2};//{'literal': 2, 'z': 8, 'op': 'literal'}
    instructions[1617] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1618] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1619] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1620] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1621] = {5'd17, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'or'}
    instructions[1622] = {5'd0, 4'd2, 4'd0, 32'd2};//{'literal': 2, 'z': 2, 'op': 'literal'}
    instructions[1623] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1624] = {5'd0, 4'd8, 4'd0, 32'd16};//{'literal': 16, 'z': 8, 'op': 'literal'}
    instructions[1625] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1626] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1627] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[1628] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[1629] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1630] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1631] = {5'd0, 4'd8, 4'd0, 32'd4};//{'literal': 4, 'z': 8, 'op': 'literal'}
    instructions[1632] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1633] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1634] = {5'd1, 4'd8, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 8, 'op': 'addl'}
    instructions[1635] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1636] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1637] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1638] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1639] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[1640] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1641] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[1642] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[1643] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1644] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1645] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1646] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1647] = {5'd16, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'shift_left'}
    instructions[1648] = {5'd0, 4'd2, 4'd0, 32'd2723};//{'literal': 2723, 'z': 2, 'op': 'literal'}
    instructions[1649] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1650] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[1651] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[1652] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1653] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1654] = {5'd0, 4'd8, 4'd0, 32'd5};//{'literal': 5, 'z': 8, 'op': 'literal'}
    instructions[1655] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1656] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1657] = {5'd1, 4'd8, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 8, 'op': 'addl'}
    instructions[1658] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1659] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1660] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1661] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1662] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[1663] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1664] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[1665] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[1666] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1667] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1668] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1669] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1670] = {5'd0, 4'd8, 4'd0, 32'd2723};//{'literal': 2723, 'z': 8, 'op': 'literal'}
    instructions[1671] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1672] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1673] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1674] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1675] = {5'd17, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'or'}
    instructions[1676] = {5'd0, 4'd2, 4'd0, 32'd2723};//{'literal': 2723, 'z': 2, 'op': 'literal'}
    instructions[1677] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1678] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[1679] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[1680] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1681] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1682] = {5'd0, 4'd8, 4'd0, 32'd7};//{'literal': 7, 'z': 8, 'op': 'literal'}
    instructions[1683] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1684] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1685] = {5'd1, 4'd8, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 8, 'op': 'addl'}
    instructions[1686] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1687] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1688] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1689] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1690] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[1691] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1692] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[1693] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[1694] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1695] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1696] = {5'd0, 4'd2, 4'd0, 32'd1};//{'literal': 1, 'z': 2, 'op': 'literal'}
    instructions[1697] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1698] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[1699] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1700] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1701] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[1702] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[1703] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1704] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1705] = {5'd0, 4'd8, 4'd0, 32'd6};//{'literal': 6, 'z': 8, 'op': 'literal'}
    instructions[1706] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1707] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1708] = {5'd1, 4'd8, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 8, 'op': 'addl'}
    instructions[1709] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1710] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1711] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1712] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1713] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[1714] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1715] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[1716] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[1717] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1718] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1719] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1720] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1721] = {5'd15, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'and'}
    instructions[1722] = {5'd0, 4'd2, 4'd0, 32'd2722};//{'literal': 2722, 'z': 2, 'op': 'literal'}
    instructions[1723] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1724] = {5'd0, 4'd8, 4'd0, 32'd2};//{'literal': 2, 'z': 8, 'op': 'literal'}
    instructions[1725] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1726] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1727] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[1728] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[1729] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1730] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1731] = {5'd0, 4'd8, 4'd0, 32'd6};//{'literal': 6, 'z': 8, 'op': 'literal'}
    instructions[1732] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1733] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1734] = {5'd1, 4'd8, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 8, 'op': 'addl'}
    instructions[1735] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1736] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1737] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1738] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1739] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[1740] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1741] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[1742] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[1743] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1744] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1745] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1746] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1747] = {5'd15, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'and'}
    instructions[1748] = {5'd0, 4'd2, 4'd0, 32'd1128};//{'literal': 1128, 'z': 2, 'op': 'literal'}
    instructions[1749] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1750] = {5'd0, 4'd8, 4'd0, 32'd4};//{'literal': 4, 'z': 8, 'op': 'literal'}
    instructions[1751] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1752] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1753] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[1754] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[1755] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1756] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1757] = {5'd0, 4'd8, 4'd0, 32'd6};//{'literal': 6, 'z': 8, 'op': 'literal'}
    instructions[1758] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1759] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1760] = {5'd1, 4'd8, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 8, 'op': 'addl'}
    instructions[1761] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1762] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1763] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1764] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1765] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[1766] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1767] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[1768] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[1769] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1770] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1771] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1772] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1773] = {5'd15, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'and'}
    instructions[1774] = {5'd0, 4'd2, 4'd0, 32'd1127};//{'literal': 1127, 'z': 2, 'op': 'literal'}
    instructions[1775] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1776] = {5'd0, 4'd8, 4'd0, 32'd8};//{'literal': 8, 'z': 8, 'op': 'literal'}
    instructions[1777] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1778] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1779] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[1780] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[1781] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1782] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1783] = {5'd0, 4'd8, 4'd0, 32'd6};//{'literal': 6, 'z': 8, 'op': 'literal'}
    instructions[1784] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1785] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1786] = {5'd1, 4'd8, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 8, 'op': 'addl'}
    instructions[1787] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1788] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1789] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1790] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1791] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[1792] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1793] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[1794] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[1795] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1796] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1797] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1798] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1799] = {5'd15, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'and'}
    instructions[1800] = {5'd0, 4'd2, 4'd0, 32'd1125};//{'literal': 1125, 'z': 2, 'op': 'literal'}
    instructions[1801] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1802] = {5'd0, 4'd8, 4'd0, 32'd16};//{'literal': 16, 'z': 8, 'op': 'literal'}
    instructions[1803] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1804] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1805] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[1806] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[1807] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1808] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1809] = {5'd0, 4'd8, 4'd0, 32'd6};//{'literal': 6, 'z': 8, 'op': 'literal'}
    instructions[1810] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1811] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1812] = {5'd1, 4'd8, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 8, 'op': 'addl'}
    instructions[1813] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1814] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1815] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1816] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1817] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[1818] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1819] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[1820] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[1821] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1822] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1823] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1824] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1825] = {5'd15, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'and'}
    instructions[1826] = {5'd0, 4'd2, 4'd0, 32'd50};//{'literal': 50, 'z': 2, 'op': 'literal'}
    instructions[1827] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1828] = {5'd0, 4'd8, 4'd0, 32'd32};//{'literal': 32, 'z': 8, 'op': 'literal'}
    instructions[1829] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1830] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1831] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[1832] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[1833] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1834] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1835] = {5'd0, 4'd8, 4'd0, 32'd6};//{'literal': 6, 'z': 8, 'op': 'literal'}
    instructions[1836] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1837] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1838] = {5'd1, 4'd8, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 8, 'op': 'addl'}
    instructions[1839] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1840] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1841] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1842] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1843] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[1844] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1845] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[1846] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[1847] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1848] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1849] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1850] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1851] = {5'd15, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'and'}
    instructions[1852] = {5'd0, 4'd2, 4'd0, 32'd52};//{'literal': 52, 'z': 2, 'op': 'literal'}
    instructions[1853] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1854] = {5'd1, 4'd8, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 8, 'op': 'addl'}
    instructions[1855] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1856] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1857] = {5'd0, 4'd2, 4'd0, 32'd2701};//{'literal': 2701, 'z': 2, 'op': 'literal'}
    instructions[1858] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1859] = {5'd1, 4'd3, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[1860] = {5'd1, 4'd4, 4'd7, 32'd0};//{'a': 7, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[1861] = {5'd12, 4'd0, 4'd6, 32'd0};//{'a': 6, 'op': 'return'}
    instructions[1862] = {5'd1, 4'd3, 4'd3, 32'd10};//{'a': 3, 'literal': 10, 'z': 3, 'op': 'addl'}
    instructions[1863] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[1864] = {5'd1, 4'd2, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1865] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1866] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[1867] = {5'd1, 4'd2, 4'd4, 32'd1};//{'a': 4, 'literal': 1, 'z': 2, 'op': 'addl'}
    instructions[1868] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1869] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[1870] = {5'd1, 4'd2, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 2, 'op': 'addl'}
    instructions[1871] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1872] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[1873] = {5'd1, 4'd2, 4'd4, 32'd3};//{'a': 4, 'literal': 3, 'z': 2, 'op': 'addl'}
    instructions[1874] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1875] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[1876] = {5'd1, 4'd2, 4'd4, 32'd4};//{'a': 4, 'literal': 4, 'z': 2, 'op': 'addl'}
    instructions[1877] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1878] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[1879] = {5'd1, 4'd2, 4'd4, 32'd5};//{'a': 4, 'literal': 5, 'z': 2, 'op': 'addl'}
    instructions[1880] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1881] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[1882] = {5'd1, 4'd2, 4'd4, 32'd6};//{'a': 4, 'literal': 6, 'z': 2, 'op': 'addl'}
    instructions[1883] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1884] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[1885] = {5'd1, 4'd2, 4'd4, 32'd7};//{'a': 4, 'literal': 7, 'z': 2, 'op': 'addl'}
    instructions[1886] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1887] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[1888] = {5'd1, 4'd2, 4'd4, 32'd8};//{'a': 4, 'literal': 8, 'z': 2, 'op': 'addl'}
    instructions[1889] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1890] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[1891] = {5'd1, 4'd2, 4'd4, 32'd9};//{'a': 4, 'literal': 9, 'z': 2, 'op': 'addl'}
    instructions[1892] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1893] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[1894] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1895] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[1896] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1897] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[1898] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[1899] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1900] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1901] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[1902] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[1903] = {5'd3, 4'd6, 4'd0, 32'd2402};//{'z': 6, 'label': 2402, 'op': 'call'}
    instructions[1904] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1905] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1906] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[1907] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1908] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[1909] = {5'd0, 4'd2, 4'd0, 32'd1092};//{'literal': 1092, 'z': 2, 'op': 'literal'}
    instructions[1910] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1911] = {5'd1, 4'd2, 4'd4, 32'd9};//{'a': 4, 'literal': 9, 'z': 2, 'op': 'addl'}
    instructions[1912] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1913] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[1914] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1915] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1916] = {5'd1, 4'd8, 4'd4, 32'd9};//{'a': 4, 'literal': 9, 'z': 8, 'op': 'addl'}
    instructions[1917] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1918] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1919] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1920] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1921] = {5'd7, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'equal'}
    instructions[1922] = {5'd6, 4'd0, 4'd8, 32'd1930};//{'a': 8, 'label': 1930, 'op': 'jmp_if_false'}
    instructions[1923] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[1924] = {5'd0, 4'd2, 4'd0, 32'd42};//{'literal': 42, 'z': 2, 'op': 'literal'}
    instructions[1925] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1926] = {5'd1, 4'd3, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[1927] = {5'd1, 4'd4, 4'd7, 32'd0};//{'a': 7, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[1928] = {5'd12, 4'd0, 4'd6, 32'd0};//{'a': 6, 'op': 'return'}
    instructions[1929] = {5'd8, 4'd0, 4'd0, 32'd1930};//{'label': 1930, 'op': 'goto'}
    instructions[1930] = {5'd0, 4'd8, 4'd0, 32'd2048};//{'literal': 2048, 'z': 8, 'op': 'literal'}
    instructions[1931] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1932] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1933] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[1934] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[1935] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1936] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1937] = {5'd0, 4'd8, 4'd0, 32'd6};//{'literal': 6, 'z': 8, 'op': 'literal'}
    instructions[1938] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1939] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[1940] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[1941] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1942] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1943] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1944] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1945] = {5'd18, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'not_equal'}
    instructions[1946] = {5'd6, 4'd0, 4'd8, 32'd1954};//{'a': 8, 'label': 1954, 'op': 'jmp_if_false'}
    instructions[1947] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[1948] = {5'd0, 4'd2, 4'd0, 32'd42};//{'literal': 42, 'z': 2, 'op': 'literal'}
    instructions[1949] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1950] = {5'd1, 4'd3, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[1951] = {5'd1, 4'd4, 4'd7, 32'd0};//{'a': 7, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[1952] = {5'd12, 4'd0, 4'd6, 32'd0};//{'a': 6, 'op': 'return'}
    instructions[1953] = {5'd8, 4'd0, 4'd0, 32'd1954};//{'label': 1954, 'op': 'goto'}
    instructions[1954] = {5'd0, 4'd8, 4'd0, 32'd49320};//{'literal': 49320, 'z': 8, 'op': 'literal'}
    instructions[1955] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1956] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1957] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[1958] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[1959] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1960] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1961] = {5'd0, 4'd8, 4'd0, 32'd15};//{'literal': 15, 'z': 8, 'op': 'literal'}
    instructions[1962] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1963] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[1964] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[1965] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1966] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1967] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1968] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1969] = {5'd18, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'not_equal'}
    instructions[1970] = {5'd6, 4'd0, 4'd8, 32'd1978};//{'a': 8, 'label': 1978, 'op': 'jmp_if_false'}
    instructions[1971] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[1972] = {5'd0, 4'd2, 4'd0, 32'd42};//{'literal': 42, 'z': 2, 'op': 'literal'}
    instructions[1973] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1974] = {5'd1, 4'd3, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[1975] = {5'd1, 4'd4, 4'd7, 32'd0};//{'a': 7, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[1976] = {5'd12, 4'd0, 4'd6, 32'd0};//{'a': 6, 'op': 'return'}
    instructions[1977] = {5'd8, 4'd0, 4'd0, 32'd1978};//{'label': 1978, 'op': 'goto'}
    instructions[1978] = {5'd0, 4'd8, 4'd0, 32'd257};//{'literal': 257, 'z': 8, 'op': 'literal'}
    instructions[1979] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1980] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1981] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[1982] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[1983] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[1984] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[1985] = {5'd0, 4'd8, 4'd0, 32'd16};//{'literal': 16, 'z': 8, 'op': 'literal'}
    instructions[1986] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1987] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[1988] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[1989] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[1990] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[1991] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1992] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[1993] = {5'd18, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'not_equal'}
    instructions[1994] = {5'd6, 4'd0, 4'd8, 32'd2002};//{'a': 8, 'label': 2002, 'op': 'jmp_if_false'}
    instructions[1995] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[1996] = {5'd0, 4'd2, 4'd0, 32'd42};//{'literal': 42, 'z': 2, 'op': 'literal'}
    instructions[1997] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[1998] = {5'd1, 4'd3, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[1999] = {5'd1, 4'd4, 4'd7, 32'd0};//{'a': 7, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[2000] = {5'd12, 4'd0, 4'd6, 32'd0};//{'a': 6, 'op': 'return'}
    instructions[2001] = {5'd8, 4'd0, 4'd0, 32'd2002};//{'label': 2002, 'op': 'goto'}
    instructions[2002] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[2003] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2004] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2005] = {5'd0, 4'd8, 4'd0, 32'd255};//{'literal': 255, 'z': 8, 'op': 'literal'}
    instructions[2006] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2007] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2008] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[2009] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[2010] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2011] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2012] = {5'd0, 4'd8, 4'd0, 32'd11};//{'literal': 11, 'z': 8, 'op': 'literal'}
    instructions[2013] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2014] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[2015] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[2016] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2017] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2018] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2019] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[2020] = {5'd15, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'and'}
    instructions[2021] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2022] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[2023] = {5'd7, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'equal'}
    instructions[2024] = {5'd6, 4'd0, 4'd8, 32'd2364};//{'a': 8, 'label': 2364, 'op': 'jmp_if_false'}
    instructions[2025] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[2026] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2027] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2028] = {5'd0, 4'd8, 4'd0, 32'd15};//{'literal': 15, 'z': 8, 'op': 'literal'}
    instructions[2029] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2030] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2031] = {5'd0, 4'd8, 4'd0, 32'd8};//{'literal': 8, 'z': 8, 'op': 'literal'}
    instructions[2032] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2033] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2034] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[2035] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[2036] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2037] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2038] = {5'd0, 4'd8, 4'd0, 32'd7};//{'literal': 7, 'z': 8, 'op': 'literal'}
    instructions[2039] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2040] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[2041] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[2042] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2043] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2044] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2045] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[2046] = {5'd14, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'unsigned_shift_right'}
    instructions[2047] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2048] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[2049] = {5'd15, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'and'}
    instructions[2050] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2051] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[2052] = {5'd16, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'shift_left'}
    instructions[2053] = {5'd1, 4'd2, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 2, 'op': 'addl'}
    instructions[2054] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[2055] = {5'd0, 4'd8, 4'd0, 32'd7};//{'literal': 7, 'z': 8, 'op': 'literal'}
    instructions[2056] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2057] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2058] = {5'd1, 4'd8, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 8, 'op': 'addl'}
    instructions[2059] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2060] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2061] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2062] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[2063] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[2064] = {5'd1, 4'd2, 4'd4, 32'd3};//{'a': 4, 'literal': 3, 'z': 2, 'op': 'addl'}
    instructions[2065] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[2066] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[2067] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[2068] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2069] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2070] = {5'd0, 4'd8, 4'd0, 32'd8};//{'literal': 8, 'z': 8, 'op': 'literal'}
    instructions[2071] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2072] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[2073] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[2074] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2075] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2076] = {5'd1, 4'd2, 4'd4, 32'd1};//{'a': 4, 'literal': 1, 'z': 2, 'op': 'addl'}
    instructions[2077] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[2078] = {5'd1, 4'd8, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 8, 'op': 'addl'}
    instructions[2079] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2080] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2081] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2082] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2083] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[2084] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2085] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2086] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[2087] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2088] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2089] = {5'd1, 4'd8, 4'd4, 32'd1};//{'a': 4, 'literal': 1, 'z': 8, 'op': 'addl'}
    instructions[2090] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2091] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2092] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2093] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[2094] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[2095] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2096] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[2097] = {5'd14, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'unsigned_shift_right'}
    instructions[2098] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2099] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[2100] = {5'd10, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'subtract'}
    instructions[2101] = {5'd1, 4'd2, 4'd4, 32'd4};//{'a': 4, 'literal': 4, 'z': 2, 'op': 'addl'}
    instructions[2102] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[2103] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[2104] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2105] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2106] = {5'd1, 4'd8, 4'd4, 32'd4};//{'a': 4, 'literal': 4, 'z': 8, 'op': 'addl'}
    instructions[2107] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2108] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2109] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2110] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2111] = {5'd1, 4'd8, 4'd4, 32'd3};//{'a': 4, 'literal': 3, 'z': 8, 'op': 'addl'}
    instructions[2112] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2113] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2114] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2115] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[2116] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[2117] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2118] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[2119] = {5'd10, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'subtract'}
    instructions[2120] = {5'd1, 4'd2, 4'd4, 32'd8};//{'a': 4, 'literal': 8, 'z': 2, 'op': 'addl'}
    instructions[2121] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[2122] = {5'd0, 4'd8, 4'd0, 32'd2048};//{'literal': 2048, 'z': 8, 'op': 'literal'}
    instructions[2123] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2124] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2125] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[2126] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[2127] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2128] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2129] = {5'd1, 4'd8, 4'd4, 32'd3};//{'a': 4, 'literal': 3, 'z': 8, 'op': 'addl'}
    instructions[2130] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2131] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2132] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2133] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[2134] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[2135] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2136] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2137] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2138] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[2139] = {5'd7, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'equal'}
    instructions[2140] = {5'd6, 4'd0, 4'd8, 32'd2357};//{'a': 8, 'label': 2357, 'op': 'jmp_if_false'}
    instructions[2141] = {5'd0, 4'd8, 4'd0, 32'd19};//{'literal': 19, 'z': 8, 'op': 'literal'}
    instructions[2142] = {5'd1, 4'd2, 4'd4, 32'd7};//{'a': 4, 'literal': 7, 'z': 2, 'op': 'addl'}
    instructions[2143] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[2144] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[2145] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2146] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[2147] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2148] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[2149] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[2150] = {5'd3, 4'd6, 4'd0, 32'd3258};//{'z': 6, 'label': 3258, 'op': 'call'}
    instructions[2151] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[2152] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2153] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[2154] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2155] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[2156] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[2157] = {5'd0, 4'd8, 4'd0, 32'd2};//{'literal': 2, 'z': 8, 'op': 'literal'}
    instructions[2158] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2159] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2160] = {5'd1, 4'd8, 4'd4, 32'd3};//{'a': 4, 'literal': 3, 'z': 8, 'op': 'addl'}
    instructions[2161] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2162] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2163] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2164] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[2165] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[2166] = {5'd1, 4'd2, 4'd4, 32'd6};//{'a': 4, 'literal': 6, 'z': 2, 'op': 'addl'}
    instructions[2167] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[2168] = {5'd1, 4'd8, 4'd4, 32'd6};//{'a': 4, 'literal': 6, 'z': 8, 'op': 'addl'}
    instructions[2169] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2170] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2171] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2172] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2173] = {5'd1, 4'd8, 4'd4, 32'd8};//{'a': 4, 'literal': 8, 'z': 8, 'op': 'addl'}
    instructions[2174] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2175] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2176] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2177] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[2178] = {5'd19, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'unsigned_greater_equal'}
    instructions[2179] = {5'd6, 4'd0, 4'd8, 32'd2267};//{'a': 8, 'label': 2267, 'op': 'jmp_if_false'}
    instructions[2180] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[2181] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[2182] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2183] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2184] = {5'd1, 4'd8, 4'd4, 32'd6};//{'a': 4, 'literal': 6, 'z': 8, 'op': 'addl'}
    instructions[2185] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2186] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2187] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2188] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[2189] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[2190] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2191] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2192] = {5'd1, 4'd2, 4'd4, 32'd5};//{'a': 4, 'literal': 5, 'z': 2, 'op': 'addl'}
    instructions[2193] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[2194] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[2195] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2196] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[2197] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2198] = {5'd1, 4'd8, 4'd4, 32'd5};//{'a': 4, 'literal': 5, 'z': 8, 'op': 'addl'}
    instructions[2199] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2200] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2201] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2202] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2203] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[2204] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[2205] = {5'd3, 4'd6, 4'd0, 32'd3268};//{'z': 6, 'label': 3268, 'op': 'call'}
    instructions[2206] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2207] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2208] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[2209] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2210] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[2211] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[2212] = {5'd1, 4'd8, 4'd4, 32'd5};//{'a': 4, 'literal': 5, 'z': 8, 'op': 'addl'}
    instructions[2213] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2214] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2215] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2216] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2217] = {5'd0, 4'd8, 4'd0, 32'd2173};//{'literal': 2173, 'z': 8, 'op': 'literal'}
    instructions[2218] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2219] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2220] = {5'd1, 4'd8, 4'd4, 32'd7};//{'a': 4, 'literal': 7, 'z': 8, 'op': 'addl'}
    instructions[2221] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2222] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2223] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2224] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[2225] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[2226] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2227] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2228] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[2229] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[2230] = {5'd1, 4'd8, 4'd4, 32'd7};//{'a': 4, 'literal': 7, 'z': 8, 'op': 'addl'}
    instructions[2231] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2232] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2233] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2234] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2235] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[2236] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2237] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2238] = {5'd1, 4'd8, 4'd4, 32'd7};//{'a': 4, 'literal': 7, 'z': 8, 'op': 'addl'}
    instructions[2239] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2240] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2241] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2242] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[2243] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[2244] = {5'd1, 4'd2, 4'd4, 32'd7};//{'a': 4, 'literal': 7, 'z': 2, 'op': 'addl'}
    instructions[2245] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[2246] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2247] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[2248] = {5'd1, 4'd8, 4'd4, 32'd6};//{'a': 4, 'literal': 6, 'z': 8, 'op': 'addl'}
    instructions[2249] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2250] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2251] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2252] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2253] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[2254] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2255] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2256] = {5'd1, 4'd8, 4'd4, 32'd6};//{'a': 4, 'literal': 6, 'z': 8, 'op': 'addl'}
    instructions[2257] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2258] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2259] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2260] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[2261] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[2262] = {5'd1, 4'd2, 4'd4, 32'd6};//{'a': 4, 'literal': 6, 'z': 2, 'op': 'addl'}
    instructions[2263] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[2264] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2265] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[2266] = {5'd8, 4'd0, 4'd0, 32'd2168};//{'label': 2168, 'op': 'goto'}
    instructions[2267] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[2268] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2269] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2270] = {5'd0, 4'd8, 4'd0, 32'd2173};//{'literal': 2173, 'z': 8, 'op': 'literal'}
    instructions[2271] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2272] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2273] = {5'd0, 4'd8, 4'd0, 32'd17};//{'literal': 17, 'z': 8, 'op': 'literal'}
    instructions[2274] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2275] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[2276] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[2277] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2278] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2279] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[2280] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[2281] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[2282] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2283] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[2284] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2285] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[2286] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[2287] = {5'd3, 4'd6, 4'd0, 32'd3357};//{'z': 6, 'label': 3357, 'op': 'call'}
    instructions[2288] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[2289] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2290] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[2291] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2292] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[2293] = {5'd0, 4'd2, 4'd0, 32'd43};//{'literal': 43, 'z': 2, 'op': 'literal'}
    instructions[2294] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2295] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2296] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2297] = {5'd0, 4'd8, 4'd0, 32'd2173};//{'literal': 2173, 'z': 8, 'op': 'literal'}
    instructions[2298] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2299] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2300] = {5'd0, 4'd8, 4'd0, 32'd18};//{'literal': 18, 'z': 8, 'op': 'literal'}
    instructions[2301] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2302] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[2303] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[2304] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2305] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2306] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[2307] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[2308] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[2309] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2310] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[2311] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2312] = {5'd0, 4'd8, 4'd0, 32'd2173};//{'literal': 2173, 'z': 8, 'op': 'literal'}
    instructions[2313] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2314] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2315] = {5'd1, 4'd8, 4'd4, 32'd1};//{'a': 4, 'literal': 1, 'z': 8, 'op': 'addl'}
    instructions[2316] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2317] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2318] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2319] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2320] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[2321] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2322] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2323] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[2324] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[2325] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2326] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2327] = {5'd0, 4'd8, 4'd0, 32'd13};//{'literal': 13, 'z': 8, 'op': 'literal'}
    instructions[2328] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2329] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[2330] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[2331] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2332] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2333] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2334] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2335] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[2336] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[2337] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2338] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2339] = {5'd0, 4'd8, 4'd0, 32'd14};//{'literal': 14, 'z': 8, 'op': 'literal'}
    instructions[2340] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2341] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[2342] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[2343] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2344] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2345] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2346] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2347] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[2348] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[2349] = {5'd3, 4'd6, 4'd0, 32'd3370};//{'z': 6, 'label': 3370, 'op': 'call'}
    instructions[2350] = {5'd1, 4'd3, 4'd3, -32'd5};//{'a': 3, 'literal': -5, 'z': 3, 'op': 'addl'}
    instructions[2351] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2352] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[2353] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2354] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[2355] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[2356] = {5'd8, 4'd0, 4'd0, 32'd2357};//{'label': 2357, 'op': 'goto'}
    instructions[2357] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[2358] = {5'd0, 4'd2, 4'd0, 32'd42};//{'literal': 42, 'z': 2, 'op': 'literal'}
    instructions[2359] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[2360] = {5'd1, 4'd3, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[2361] = {5'd1, 4'd4, 4'd7, 32'd0};//{'a': 7, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[2362] = {5'd12, 4'd0, 4'd6, 32'd0};//{'a': 6, 'op': 'return'}
    instructions[2363] = {5'd8, 4'd0, 4'd0, 32'd2364};//{'label': 2364, 'op': 'goto'}
    instructions[2364] = {5'd0, 4'd8, 4'd0, 32'd6};//{'literal': 6, 'z': 8, 'op': 'literal'}
    instructions[2365] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2366] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2367] = {5'd0, 4'd8, 4'd0, 32'd255};//{'literal': 255, 'z': 8, 'op': 'literal'}
    instructions[2368] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2369] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2370] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[2371] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[2372] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2373] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2374] = {5'd0, 4'd8, 4'd0, 32'd11};//{'literal': 11, 'z': 8, 'op': 'literal'}
    instructions[2375] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2376] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[2377] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[2378] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2379] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2380] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2381] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[2382] = {5'd15, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'and'}
    instructions[2383] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2384] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[2385] = {5'd18, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'not_equal'}
    instructions[2386] = {5'd6, 4'd0, 4'd8, 32'd2394};//{'a': 8, 'label': 2394, 'op': 'jmp_if_false'}
    instructions[2387] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[2388] = {5'd0, 4'd2, 4'd0, 32'd42};//{'literal': 42, 'z': 2, 'op': 'literal'}
    instructions[2389] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[2390] = {5'd1, 4'd3, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[2391] = {5'd1, 4'd4, 4'd7, 32'd0};//{'a': 7, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[2392] = {5'd12, 4'd0, 4'd6, 32'd0};//{'a': 6, 'op': 'return'}
    instructions[2393] = {5'd8, 4'd0, 4'd0, 32'd2394};//{'label': 2394, 'op': 'goto'}
    instructions[2394] = {5'd1, 4'd8, 4'd4, 32'd9};//{'a': 4, 'literal': 9, 'z': 8, 'op': 'addl'}
    instructions[2395] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2396] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2397] = {5'd0, 4'd2, 4'd0, 32'd42};//{'literal': 42, 'z': 2, 'op': 'literal'}
    instructions[2398] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[2399] = {5'd1, 4'd3, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[2400] = {5'd1, 4'd4, 4'd7, 32'd0};//{'a': 7, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[2401] = {5'd12, 4'd0, 4'd6, 32'd0};//{'a': 6, 'op': 'return'}
    instructions[2402] = {5'd1, 4'd3, 4'd3, 32'd3};//{'a': 3, 'literal': 3, 'z': 3, 'op': 'addl'}
    instructions[2403] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[2404] = {5'd1, 4'd2, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2405] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[2406] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[2407] = {5'd1, 4'd2, 4'd4, 32'd1};//{'a': 4, 'literal': 1, 'z': 2, 'op': 'addl'}
    instructions[2408] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[2409] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[2410] = {5'd1, 4'd2, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 2, 'op': 'addl'}
    instructions[2411] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[2412] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[2413] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2414] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2415] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[2416] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2417] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[2418] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2419] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[2420] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[2421] = {5'd3, 4'd6, 4'd0, 32'd3006};//{'z': 6, 'label': 3006, 'op': 'call'}
    instructions[2422] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[2423] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2424] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[2425] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2426] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[2427] = {5'd0, 4'd2, 4'd0, 32'd0};//{'literal': 0, 'z': 2, 'op': 'literal'}
    instructions[2428] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2429] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2430] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[2431] = {5'd7, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'equal'}
    instructions[2432] = {5'd6, 4'd0, 4'd8, 32'd2440};//{'a': 8, 'label': 2440, 'op': 'jmp_if_false'}
    instructions[2433] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[2434] = {5'd0, 4'd2, 4'd0, 32'd1092};//{'literal': 1092, 'z': 2, 'op': 'literal'}
    instructions[2435] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[2436] = {5'd1, 4'd3, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[2437] = {5'd1, 4'd4, 4'd7, 32'd0};//{'a': 7, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[2438] = {5'd12, 4'd0, 4'd6, 32'd0};//{'a': 6, 'op': 'return'}
    instructions[2439] = {5'd8, 4'd0, 4'd0, 32'd2440};//{'label': 2440, 'op': 'goto'}
    instructions[2440] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[2441] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2442] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[2443] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2444] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[2445] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[2446] = {5'd3, 4'd6, 4'd0, 32'd3016};//{'z': 6, 'label': 3016, 'op': 'call'}
    instructions[2447] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[2448] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2449] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[2450] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2451] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[2452] = {5'd0, 4'd2, 4'd0, 32'd1081};//{'literal': 1081, 'z': 2, 'op': 'literal'}
    instructions[2453] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2454] = {5'd1, 4'd2, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2455] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[2456] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[2457] = {5'd1, 4'd2, 4'd4, 32'd1};//{'a': 4, 'literal': 1, 'z': 2, 'op': 'addl'}
    instructions[2458] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[2459] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[2460] = {5'd1, 4'd2, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 2, 'op': 'addl'}
    instructions[2461] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[2462] = {5'd1, 4'd8, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 8, 'op': 'addl'}
    instructions[2463] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2464] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2465] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2466] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2467] = {5'd1, 4'd8, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 8, 'op': 'addl'}
    instructions[2468] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2469] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2470] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2471] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[2472] = {5'd20, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'unsigned_greater'}
    instructions[2473] = {5'd6, 4'd0, 4'd8, 32'd2534};//{'a': 8, 'label': 2534, 'op': 'jmp_if_false'}
    instructions[2474] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[2475] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2476] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[2477] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2478] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[2479] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[2480] = {5'd3, 4'd6, 4'd0, 32'd3016};//{'z': 6, 'label': 3016, 'op': 'call'}
    instructions[2481] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[2482] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2483] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[2484] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2485] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[2486] = {5'd0, 4'd2, 4'd0, 32'd1081};//{'literal': 1081, 'z': 2, 'op': 'literal'}
    instructions[2487] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2488] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2489] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2490] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[2491] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[2492] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2493] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2494] = {5'd1, 4'd8, 4'd4, 32'd1};//{'a': 4, 'literal': 1, 'z': 8, 'op': 'addl'}
    instructions[2495] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2496] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2497] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2498] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[2499] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[2500] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2501] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2502] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[2503] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[2504] = {5'd1, 4'd8, 4'd4, 32'd1};//{'a': 4, 'literal': 1, 'z': 8, 'op': 'addl'}
    instructions[2505] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2506] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2507] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2508] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2509] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[2510] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2511] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2512] = {5'd1, 4'd8, 4'd4, 32'd1};//{'a': 4, 'literal': 1, 'z': 8, 'op': 'addl'}
    instructions[2513] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2514] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2515] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2516] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[2517] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[2518] = {5'd1, 4'd2, 4'd4, 32'd1};//{'a': 4, 'literal': 1, 'z': 2, 'op': 'addl'}
    instructions[2519] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[2520] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2521] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[2522] = {5'd0, 4'd8, 4'd0, 32'd2};//{'literal': 2, 'z': 8, 'op': 'literal'}
    instructions[2523] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2524] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2525] = {5'd1, 4'd8, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 8, 'op': 'addl'}
    instructions[2526] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2527] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2528] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2529] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[2530] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[2531] = {5'd1, 4'd2, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 2, 'op': 'addl'}
    instructions[2532] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[2533] = {5'd8, 4'd0, 4'd0, 32'd2462};//{'label': 2462, 'op': 'goto'}
    instructions[2534] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[2535] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2536] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2537] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[2538] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[2539] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2540] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2541] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[2542] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2543] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[2544] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[2545] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2546] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2547] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2548] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[2549] = {5'd18, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'not_equal'}
    instructions[2550] = {5'd6, 4'd0, 4'd8, 32'd2567};//{'a': 8, 'label': 2567, 'op': 'jmp_if_false'}
    instructions[2551] = {5'd0, 4'd8, 4'd0, 32'd65535};//{'literal': 65535, 'z': 8, 'op': 'literal'}
    instructions[2552] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2553] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2554] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[2555] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[2556] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2557] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2558] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[2559] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2560] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[2561] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[2562] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2563] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2564] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2565] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[2566] = {5'd18, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'not_equal'}
    instructions[2567] = {5'd6, 4'd0, 4'd8, 32'd2575};//{'a': 8, 'label': 2575, 'op': 'jmp_if_false'}
    instructions[2568] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[2569] = {5'd0, 4'd2, 4'd0, 32'd1092};//{'literal': 1092, 'z': 2, 'op': 'literal'}
    instructions[2570] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[2571] = {5'd1, 4'd3, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[2572] = {5'd1, 4'd4, 4'd7, 32'd0};//{'a': 7, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[2573] = {5'd12, 4'd0, 4'd6, 32'd0};//{'a': 6, 'op': 'return'}
    instructions[2574] = {5'd8, 4'd0, 4'd0, 32'd2575};//{'label': 2575, 'op': 'goto'}
    instructions[2575] = {5'd0, 4'd8, 4'd0, 32'd515};//{'literal': 515, 'z': 8, 'op': 'literal'}
    instructions[2576] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2577] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2578] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[2579] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[2580] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2581] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2582] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[2583] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2584] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[2585] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[2586] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2587] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2588] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2589] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[2590] = {5'd18, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'not_equal'}
    instructions[2591] = {5'd6, 4'd0, 4'd8, 32'd2608};//{'a': 8, 'label': 2608, 'op': 'jmp_if_false'}
    instructions[2592] = {5'd0, 4'd8, 4'd0, 32'd65535};//{'literal': 65535, 'z': 8, 'op': 'literal'}
    instructions[2593] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2594] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2595] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[2596] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[2597] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2598] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2599] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[2600] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2601] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[2602] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[2603] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2604] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2605] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2606] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[2607] = {5'd18, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'not_equal'}
    instructions[2608] = {5'd6, 4'd0, 4'd8, 32'd2616};//{'a': 8, 'label': 2616, 'op': 'jmp_if_false'}
    instructions[2609] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[2610] = {5'd0, 4'd2, 4'd0, 32'd1092};//{'literal': 1092, 'z': 2, 'op': 'literal'}
    instructions[2611] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[2612] = {5'd1, 4'd3, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[2613] = {5'd1, 4'd4, 4'd7, 32'd0};//{'a': 7, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[2614] = {5'd12, 4'd0, 4'd6, 32'd0};//{'a': 6, 'op': 'return'}
    instructions[2615] = {5'd8, 4'd0, 4'd0, 32'd2616};//{'label': 2616, 'op': 'goto'}
    instructions[2616] = {5'd0, 4'd8, 4'd0, 32'd1029};//{'literal': 1029, 'z': 8, 'op': 'literal'}
    instructions[2617] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2618] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2619] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[2620] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[2621] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2622] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2623] = {5'd0, 4'd8, 4'd0, 32'd2};//{'literal': 2, 'z': 8, 'op': 'literal'}
    instructions[2624] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2625] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[2626] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[2627] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2628] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2629] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2630] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[2631] = {5'd18, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'not_equal'}
    instructions[2632] = {5'd6, 4'd0, 4'd8, 32'd2649};//{'a': 8, 'label': 2649, 'op': 'jmp_if_false'}
    instructions[2633] = {5'd0, 4'd8, 4'd0, 32'd65535};//{'literal': 65535, 'z': 8, 'op': 'literal'}
    instructions[2634] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2635] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2636] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[2637] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[2638] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2639] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2640] = {5'd0, 4'd8, 4'd0, 32'd2};//{'literal': 2, 'z': 8, 'op': 'literal'}
    instructions[2641] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2642] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[2643] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[2644] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2645] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2646] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2647] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[2648] = {5'd18, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'not_equal'}
    instructions[2649] = {5'd6, 4'd0, 4'd8, 32'd2657};//{'a': 8, 'label': 2657, 'op': 'jmp_if_false'}
    instructions[2650] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[2651] = {5'd0, 4'd2, 4'd0, 32'd1092};//{'literal': 1092, 'z': 2, 'op': 'literal'}
    instructions[2652] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[2653] = {5'd1, 4'd3, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[2654] = {5'd1, 4'd4, 4'd7, 32'd0};//{'a': 7, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[2655] = {5'd12, 4'd0, 4'd6, 32'd0};//{'a': 6, 'op': 'return'}
    instructions[2656] = {5'd8, 4'd0, 4'd0, 32'd2657};//{'label': 2657, 'op': 'goto'}
    instructions[2657] = {5'd0, 4'd8, 4'd0, 32'd2054};//{'literal': 2054, 'z': 8, 'op': 'literal'}
    instructions[2658] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2659] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2660] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[2661] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[2662] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2663] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2664] = {5'd0, 4'd8, 4'd0, 32'd6};//{'literal': 6, 'z': 8, 'op': 'literal'}
    instructions[2665] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2666] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[2667] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[2668] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2669] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2670] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2671] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[2672] = {5'd7, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'equal'}
    instructions[2673] = {5'd6, 4'd0, 4'd8, 32'd2998};//{'a': 8, 'label': 2998, 'op': 'jmp_if_false'}
    instructions[2674] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[2675] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2676] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2677] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[2678] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[2679] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2680] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2681] = {5'd0, 4'd8, 4'd0, 32'd10};//{'literal': 10, 'z': 8, 'op': 'literal'}
    instructions[2682] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2683] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[2684] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[2685] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2686] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2687] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2688] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[2689] = {5'd7, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'equal'}
    instructions[2690] = {5'd6, 4'd0, 4'd8, 32'd2991};//{'a': 8, 'label': 2991, 'op': 'jmp_if_false'}
    instructions[2691] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[2692] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2693] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2694] = {5'd0, 4'd8, 4'd0, 32'd2173};//{'literal': 2173, 'z': 8, 'op': 'literal'}
    instructions[2695] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2696] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2697] = {5'd0, 4'd8, 4'd0, 32'd7};//{'literal': 7, 'z': 8, 'op': 'literal'}
    instructions[2698] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2699] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[2700] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[2701] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2702] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2703] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[2704] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[2705] = {5'd0, 4'd8, 4'd0, 32'd2048};//{'literal': 2048, 'z': 8, 'op': 'literal'}
    instructions[2706] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2707] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2708] = {5'd0, 4'd8, 4'd0, 32'd2173};//{'literal': 2173, 'z': 8, 'op': 'literal'}
    instructions[2709] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2710] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2711] = {5'd0, 4'd8, 4'd0, 32'd8};//{'literal': 8, 'z': 8, 'op': 'literal'}
    instructions[2712] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2713] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[2714] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[2715] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2716] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2717] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[2718] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[2719] = {5'd0, 4'd8, 4'd0, 32'd1540};//{'literal': 1540, 'z': 8, 'op': 'literal'}
    instructions[2720] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2721] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2722] = {5'd0, 4'd8, 4'd0, 32'd2173};//{'literal': 2173, 'z': 8, 'op': 'literal'}
    instructions[2723] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2724] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2725] = {5'd0, 4'd8, 4'd0, 32'd9};//{'literal': 9, 'z': 8, 'op': 'literal'}
    instructions[2726] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2727] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[2728] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[2729] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2730] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2731] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[2732] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[2733] = {5'd0, 4'd8, 4'd0, 32'd2};//{'literal': 2, 'z': 8, 'op': 'literal'}
    instructions[2734] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2735] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2736] = {5'd0, 4'd8, 4'd0, 32'd2173};//{'literal': 2173, 'z': 8, 'op': 'literal'}
    instructions[2737] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2738] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2739] = {5'd0, 4'd8, 4'd0, 32'd10};//{'literal': 10, 'z': 8, 'op': 'literal'}
    instructions[2740] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2741] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[2742] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[2743] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2744] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2745] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[2746] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[2747] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[2748] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2749] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2750] = {5'd0, 4'd8, 4'd0, 32'd2173};//{'literal': 2173, 'z': 8, 'op': 'literal'}
    instructions[2751] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2752] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2753] = {5'd0, 4'd8, 4'd0, 32'd11};//{'literal': 11, 'z': 8, 'op': 'literal'}
    instructions[2754] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2755] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[2756] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[2757] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2758] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2759] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[2760] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[2761] = {5'd0, 4'd8, 4'd0, 32'd515};//{'literal': 515, 'z': 8, 'op': 'literal'}
    instructions[2762] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2763] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2764] = {5'd0, 4'd8, 4'd0, 32'd2173};//{'literal': 2173, 'z': 8, 'op': 'literal'}
    instructions[2765] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2766] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2767] = {5'd0, 4'd8, 4'd0, 32'd12};//{'literal': 12, 'z': 8, 'op': 'literal'}
    instructions[2768] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2769] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[2770] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[2771] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2772] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2773] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[2774] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[2775] = {5'd0, 4'd8, 4'd0, 32'd1029};//{'literal': 1029, 'z': 8, 'op': 'literal'}
    instructions[2776] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2777] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2778] = {5'd0, 4'd8, 4'd0, 32'd2173};//{'literal': 2173, 'z': 8, 'op': 'literal'}
    instructions[2779] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2780] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2781] = {5'd0, 4'd8, 4'd0, 32'd13};//{'literal': 13, 'z': 8, 'op': 'literal'}
    instructions[2782] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2783] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[2784] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[2785] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2786] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2787] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[2788] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[2789] = {5'd0, 4'd8, 4'd0, 32'd49320};//{'literal': 49320, 'z': 8, 'op': 'literal'}
    instructions[2790] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2791] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2792] = {5'd0, 4'd8, 4'd0, 32'd2173};//{'literal': 2173, 'z': 8, 'op': 'literal'}
    instructions[2793] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2794] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2795] = {5'd0, 4'd8, 4'd0, 32'd14};//{'literal': 14, 'z': 8, 'op': 'literal'}
    instructions[2796] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2797] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[2798] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[2799] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2800] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2801] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[2802] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[2803] = {5'd0, 4'd8, 4'd0, 32'd257};//{'literal': 257, 'z': 8, 'op': 'literal'}
    instructions[2804] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2805] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2806] = {5'd0, 4'd8, 4'd0, 32'd2173};//{'literal': 2173, 'z': 8, 'op': 'literal'}
    instructions[2807] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2808] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2809] = {5'd0, 4'd8, 4'd0, 32'd15};//{'literal': 15, 'z': 8, 'op': 'literal'}
    instructions[2810] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2811] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[2812] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[2813] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2814] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2815] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[2816] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[2817] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[2818] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[2819] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2820] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2821] = {5'd0, 4'd8, 4'd0, 32'd11};//{'literal': 11, 'z': 8, 'op': 'literal'}
    instructions[2822] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2823] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[2824] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[2825] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2826] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2827] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2828] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2829] = {5'd0, 4'd8, 4'd0, 32'd2173};//{'literal': 2173, 'z': 8, 'op': 'literal'}
    instructions[2830] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2831] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2832] = {5'd0, 4'd8, 4'd0, 32'd16};//{'literal': 16, 'z': 8, 'op': 'literal'}
    instructions[2833] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2834] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[2835] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[2836] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2837] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2838] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[2839] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[2840] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[2841] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[2842] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2843] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2844] = {5'd0, 4'd8, 4'd0, 32'd12};//{'literal': 12, 'z': 8, 'op': 'literal'}
    instructions[2845] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2846] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[2847] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[2848] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2849] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2850] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2851] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2852] = {5'd0, 4'd8, 4'd0, 32'd2173};//{'literal': 2173, 'z': 8, 'op': 'literal'}
    instructions[2853] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2854] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2855] = {5'd0, 4'd8, 4'd0, 32'd17};//{'literal': 17, 'z': 8, 'op': 'literal'}
    instructions[2856] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2857] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[2858] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[2859] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2860] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2861] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[2862] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[2863] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[2864] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[2865] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2866] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2867] = {5'd0, 4'd8, 4'd0, 32'd13};//{'literal': 13, 'z': 8, 'op': 'literal'}
    instructions[2868] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2869] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[2870] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[2871] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2872] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2873] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2874] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2875] = {5'd0, 4'd8, 4'd0, 32'd2173};//{'literal': 2173, 'z': 8, 'op': 'literal'}
    instructions[2876] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2877] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2878] = {5'd0, 4'd8, 4'd0, 32'd18};//{'literal': 18, 'z': 8, 'op': 'literal'}
    instructions[2879] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2880] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[2881] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[2882] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2883] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2884] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[2885] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[2886] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[2887] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[2888] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2889] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2890] = {5'd0, 4'd8, 4'd0, 32'd14};//{'literal': 14, 'z': 8, 'op': 'literal'}
    instructions[2891] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2892] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[2893] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[2894] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2895] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2896] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2897] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2898] = {5'd0, 4'd8, 4'd0, 32'd2173};//{'literal': 2173, 'z': 8, 'op': 'literal'}
    instructions[2899] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2900] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2901] = {5'd0, 4'd8, 4'd0, 32'd19};//{'literal': 19, 'z': 8, 'op': 'literal'}
    instructions[2902] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2903] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[2904] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[2905] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2906] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2907] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[2908] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[2909] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[2910] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[2911] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2912] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2913] = {5'd0, 4'd8, 4'd0, 32'd15};//{'literal': 15, 'z': 8, 'op': 'literal'}
    instructions[2914] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2915] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[2916] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[2917] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2918] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2919] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2920] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2921] = {5'd0, 4'd8, 4'd0, 32'd2173};//{'literal': 2173, 'z': 8, 'op': 'literal'}
    instructions[2922] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2923] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2924] = {5'd0, 4'd8, 4'd0, 32'd20};//{'literal': 20, 'z': 8, 'op': 'literal'}
    instructions[2925] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2926] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[2927] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[2928] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2929] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2930] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[2931] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[2932] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[2933] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2934] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[2935] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2936] = {5'd0, 4'd8, 4'd0, 32'd2173};//{'literal': 2173, 'z': 8, 'op': 'literal'}
    instructions[2937] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2938] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2939] = {5'd0, 4'd8, 4'd0, 32'd64};//{'literal': 64, 'z': 8, 'op': 'literal'}
    instructions[2940] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2941] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2942] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[2943] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[2944] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2945] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2946] = {5'd0, 4'd8, 4'd0, 32'd11};//{'literal': 11, 'z': 8, 'op': 'literal'}
    instructions[2947] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2948] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[2949] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[2950] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2951] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2952] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2953] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2954] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[2955] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[2956] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2957] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2958] = {5'd0, 4'd8, 4'd0, 32'd12};//{'literal': 12, 'z': 8, 'op': 'literal'}
    instructions[2959] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2960] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[2961] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[2962] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2963] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2964] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2965] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2966] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[2967] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[2968] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2969] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2970] = {5'd0, 4'd8, 4'd0, 32'd13};//{'literal': 13, 'z': 8, 'op': 'literal'}
    instructions[2971] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2972] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[2973] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[2974] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[2975] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[2976] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2977] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2978] = {5'd0, 4'd8, 4'd0, 32'd2054};//{'literal': 2054, 'z': 8, 'op': 'literal'}
    instructions[2979] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[2980] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[2981] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[2982] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[2983] = {5'd3, 4'd6, 4'd0, 32'd3026};//{'z': 6, 'label': 3026, 'op': 'call'}
    instructions[2984] = {5'd1, 4'd3, 4'd3, -32'd6};//{'a': 3, 'literal': -6, 'z': 3, 'op': 'addl'}
    instructions[2985] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2986] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[2987] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[2988] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[2989] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[2990] = {5'd8, 4'd0, 4'd0, 32'd2991};//{'label': 2991, 'op': 'goto'}
    instructions[2991] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[2992] = {5'd0, 4'd2, 4'd0, 32'd1092};//{'literal': 1092, 'z': 2, 'op': 'literal'}
    instructions[2993] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[2994] = {5'd1, 4'd3, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[2995] = {5'd1, 4'd4, 4'd7, 32'd0};//{'a': 7, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[2996] = {5'd12, 4'd0, 4'd6, 32'd0};//{'a': 6, 'op': 'return'}
    instructions[2997] = {5'd8, 4'd0, 4'd0, 32'd2998};//{'label': 2998, 'op': 'goto'}
    instructions[2998] = {5'd1, 4'd8, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 8, 'op': 'addl'}
    instructions[2999] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3000] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3001] = {5'd0, 4'd2, 4'd0, 32'd1092};//{'literal': 1092, 'z': 2, 'op': 'literal'}
    instructions[3002] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3003] = {5'd1, 4'd3, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[3004] = {5'd1, 4'd4, 4'd7, 32'd0};//{'a': 7, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[3005] = {5'd12, 4'd0, 4'd6, 32'd0};//{'a': 6, 'op': 'return'}
    instructions[3006] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[3007] = {5'd0, 4'd8, 4'd0, 32'd2725};//{'literal': 2725, 'z': 8, 'op': 'literal'}
    instructions[3008] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3009] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3010] = {5'd21, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'ready'}
    instructions[3011] = {5'd0, 4'd2, 4'd0, 32'd0};//{'literal': 0, 'z': 2, 'op': 'literal'}
    instructions[3012] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3013] = {5'd1, 4'd3, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[3014] = {5'd1, 4'd4, 4'd7, 32'd0};//{'a': 7, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[3015] = {5'd12, 4'd0, 4'd6, 32'd0};//{'a': 6, 'op': 'return'}
    instructions[3016] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[3017] = {5'd0, 4'd8, 4'd0, 32'd2725};//{'literal': 2725, 'z': 8, 'op': 'literal'}
    instructions[3018] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3019] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3020] = {5'd22, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'read'}
    instructions[3021] = {5'd0, 4'd2, 4'd0, 32'd1081};//{'literal': 1081, 'z': 2, 'op': 'literal'}
    instructions[3022] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3023] = {5'd1, 4'd3, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[3024] = {5'd1, 4'd4, 4'd7, 32'd0};//{'a': 7, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[3025] = {5'd12, 4'd0, 4'd6, 32'd0};//{'a': 6, 'op': 'return'}
    instructions[3026] = {5'd1, 4'd3, 4'd3, 32'd2};//{'a': 3, 'literal': 2, 'z': 3, 'op': 'addl'}
    instructions[3027] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[3028] = {5'd1, 4'd2, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3029] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3030] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[3031] = {5'd1, 4'd2, 4'd4, 32'd1};//{'a': 4, 'literal': 1, 'z': 2, 'op': 'addl'}
    instructions[3032] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3033] = {5'd1, 4'd8, 4'd4, -32'd4};//{'a': 4, 'literal': -4, 'z': 8, 'op': 'addl'}
    instructions[3034] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3035] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3036] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3037] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3038] = {5'd1, 4'd8, 4'd4, -32'd6};//{'a': 4, 'literal': -6, 'z': 8, 'op': 'addl'}
    instructions[3039] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[3040] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3041] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3042] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[3043] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3044] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[3045] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[3046] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3047] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3048] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[3049] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3050] = {5'd1, 4'd8, 4'd4, -32'd3};//{'a': 4, 'literal': -3, 'z': 8, 'op': 'addl'}
    instructions[3051] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3052] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3053] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3054] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3055] = {5'd1, 4'd8, 4'd4, -32'd6};//{'a': 4, 'literal': -6, 'z': 8, 'op': 'addl'}
    instructions[3056] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[3057] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3058] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3059] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[3060] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3061] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[3062] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[3063] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3064] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3065] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[3066] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3067] = {5'd1, 4'd8, 4'd4, -32'd2};//{'a': 4, 'literal': -2, 'z': 8, 'op': 'addl'}
    instructions[3068] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3069] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3070] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3071] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3072] = {5'd1, 4'd8, 4'd4, -32'd6};//{'a': 4, 'literal': -6, 'z': 8, 'op': 'addl'}
    instructions[3073] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[3074] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3075] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3076] = {5'd0, 4'd8, 4'd0, 32'd2};//{'literal': 2, 'z': 8, 'op': 'literal'}
    instructions[3077] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3078] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[3079] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[3080] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3081] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3082] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[3083] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3084] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[3085] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3086] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3087] = {5'd1, 4'd8, 4'd4, -32'd6};//{'a': 4, 'literal': -6, 'z': 8, 'op': 'addl'}
    instructions[3088] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[3089] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3090] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3091] = {5'd0, 4'd8, 4'd0, 32'd3};//{'literal': 3, 'z': 8, 'op': 'literal'}
    instructions[3092] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3093] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[3094] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[3095] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3096] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3097] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[3098] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3099] = {5'd0, 4'd8, 4'd0, 32'd515};//{'literal': 515, 'z': 8, 'op': 'literal'}
    instructions[3100] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3101] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3102] = {5'd1, 4'd8, 4'd4, -32'd6};//{'a': 4, 'literal': -6, 'z': 8, 'op': 'addl'}
    instructions[3103] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[3104] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3105] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3106] = {5'd0, 4'd8, 4'd0, 32'd4};//{'literal': 4, 'z': 8, 'op': 'literal'}
    instructions[3107] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3108] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[3109] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[3110] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3111] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3112] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[3113] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3114] = {5'd0, 4'd8, 4'd0, 32'd1029};//{'literal': 1029, 'z': 8, 'op': 'literal'}
    instructions[3115] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3116] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3117] = {5'd1, 4'd8, 4'd4, -32'd6};//{'a': 4, 'literal': -6, 'z': 8, 'op': 'addl'}
    instructions[3118] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[3119] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3120] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3121] = {5'd0, 4'd8, 4'd0, 32'd5};//{'literal': 5, 'z': 8, 'op': 'literal'}
    instructions[3122] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3123] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[3124] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[3125] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3126] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3127] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[3128] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3129] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[3130] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3131] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3132] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3133] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3134] = {5'd1, 4'd8, 4'd4, -32'd6};//{'a': 4, 'literal': -6, 'z': 8, 'op': 'addl'}
    instructions[3135] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[3136] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3137] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3138] = {5'd0, 4'd8, 4'd0, 32'd6};//{'literal': 6, 'z': 8, 'op': 'literal'}
    instructions[3139] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3140] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[3141] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[3142] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3143] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3144] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[3145] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3146] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[3147] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3148] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[3149] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3150] = {5'd1, 4'd8, 4'd4, -32'd5};//{'a': 4, 'literal': -5, 'z': 8, 'op': 'addl'}
    instructions[3151] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3152] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3153] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3154] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3155] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[3156] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[3157] = {5'd3, 4'd6, 4'd0, 32'd3242};//{'z': 6, 'label': 3242, 'op': 'call'}
    instructions[3158] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3159] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3160] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[3161] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3162] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[3163] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[3164] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[3165] = {5'd1, 4'd2, 4'd4, 32'd1};//{'a': 4, 'literal': 1, 'z': 2, 'op': 'addl'}
    instructions[3166] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3167] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[3168] = {5'd1, 4'd2, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3169] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3170] = {5'd1, 4'd8, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 8, 'op': 'addl'}
    instructions[3171] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3172] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3173] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3174] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3175] = {5'd1, 4'd8, 4'd4, -32'd5};//{'a': 4, 'literal': -5, 'z': 8, 'op': 'addl'}
    instructions[3176] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3177] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3178] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3179] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[3180] = {5'd20, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'unsigned_greater'}
    instructions[3181] = {5'd6, 4'd0, 4'd8, 32'd3239};//{'a': 8, 'label': 3239, 'op': 'jmp_if_false'}
    instructions[3182] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[3183] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3184] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[3185] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3186] = {5'd1, 4'd8, 4'd4, -32'd6};//{'a': 4, 'literal': -6, 'z': 8, 'op': 'addl'}
    instructions[3187] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[3188] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3189] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3190] = {5'd1, 4'd8, 4'd4, 32'd1};//{'a': 4, 'literal': 1, 'z': 8, 'op': 'addl'}
    instructions[3191] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3192] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3193] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3194] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[3195] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[3196] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3197] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3198] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3199] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3200] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[3201] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[3202] = {5'd3, 4'd6, 4'd0, 32'd3242};//{'z': 6, 'label': 3242, 'op': 'call'}
    instructions[3203] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3204] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3205] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[3206] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3207] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[3208] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[3209] = {5'd1, 4'd8, 4'd4, 32'd1};//{'a': 4, 'literal': 1, 'z': 8, 'op': 'addl'}
    instructions[3210] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3211] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3212] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3213] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3214] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[3215] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3216] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3217] = {5'd1, 4'd8, 4'd4, 32'd1};//{'a': 4, 'literal': 1, 'z': 8, 'op': 'addl'}
    instructions[3218] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3219] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3220] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3221] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[3222] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[3223] = {5'd1, 4'd2, 4'd4, 32'd1};//{'a': 4, 'literal': 1, 'z': 2, 'op': 'addl'}
    instructions[3224] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3225] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3226] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[3227] = {5'd0, 4'd8, 4'd0, 32'd2};//{'literal': 2, 'z': 8, 'op': 'literal'}
    instructions[3228] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3229] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3230] = {5'd1, 4'd8, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 8, 'op': 'addl'}
    instructions[3231] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3232] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3233] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3234] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[3235] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[3236] = {5'd1, 4'd2, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3237] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3238] = {5'd8, 4'd0, 4'd0, 32'd3170};//{'label': 3170, 'op': 'goto'}
    instructions[3239] = {5'd1, 4'd3, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[3240] = {5'd1, 4'd4, 4'd7, 32'd0};//{'a': 7, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[3241] = {5'd12, 4'd0, 4'd6, 32'd0};//{'a': 6, 'op': 'return'}
    instructions[3242] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[3243] = {5'd0, 4'd8, 4'd0, 32'd36};//{'literal': 36, 'z': 8, 'op': 'literal'}
    instructions[3244] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3245] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3246] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3247] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3248] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[3249] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3250] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3251] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3252] = {5'd5, 4'd0, 4'd3, 32'd0};//{'a': 3, 'z': 0, 'op': 'load'}
    instructions[3253] = {5'd13, 4'd0, 4'd0, 32'd8};//{'a': 0, 'b': 8, 'op': 'write'}
    instructions[3254] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[3255] = {5'd1, 4'd3, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[3256] = {5'd1, 4'd4, 4'd7, 32'd0};//{'a': 7, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[3257] = {5'd12, 4'd0, 4'd6, 32'd0};//{'a': 6, 'op': 'return'}
    instructions[3258] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[3259] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[3260] = {5'd23, 4'd9, 4'd8, 32'd0};//{'a': 8, 'z': 9, 'op': 'int_to_long'}
    instructions[3261] = {5'd0, 4'd2, 4'd0, 32'd38};//{'literal': 38, 'z': 2, 'op': 'literal'}
    instructions[3262] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3263] = {5'd1, 4'd2, 4'd2, 32'd1};//{'a': 2, 'literal': 1, 'z': 2, 'op': 'addl'}
    instructions[3264] = {5'd2, 4'd0, 4'd2, 32'd9};//{'a': 2, 'b': 9, 'op': 'store'}
    instructions[3265] = {5'd1, 4'd3, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[3266] = {5'd1, 4'd4, 4'd7, 32'd0};//{'a': 7, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[3267] = {5'd12, 4'd0, 4'd6, 32'd0};//{'a': 6, 'op': 'return'}
    instructions[3268] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[3269] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[3270] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3271] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3272] = {5'd0, 4'd9, 4'd0, 32'd0};//{'literal': 0, 'z': 9, 'op': 'literal'}
    instructions[3273] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3274] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3275] = {5'd2, 4'd0, 4'd3, 32'd9};//{'a': 3, 'comment': 'push', 'b': 9, 'op': 'store'}
    instructions[3276] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3277] = {5'd0, 4'd8, 4'd0, 32'd38};//{'literal': 38, 'z': 8, 'op': 'literal'}
    instructions[3278] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3279] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3280] = {5'd1, 4'd2, 4'd2, 32'd1};//{'a': 2, 'literal': 1, 'z': 2, 'op': 'addl'}
    instructions[3281] = {5'd5, 4'd9, 4'd2, 32'd0};//{'a': 2, 'z': 9, 'op': 'load'}
    instructions[3282] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3283] = {5'd5, 4'd11, 4'd3, 32'd0};//{'a': 3, 'z': 11, 'op': 'load'}
    instructions[3284] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3285] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[3286] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[3287] = {5'd24, 4'd9, 4'd9, 32'd11};//{'a': 9, 'z': 9, 'b': 11, 'op': 'add_with_carry'}
    instructions[3288] = {5'd0, 4'd2, 4'd0, 32'd38};//{'literal': 38, 'z': 2, 'op': 'literal'}
    instructions[3289] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3290] = {5'd1, 4'd2, 4'd2, 32'd1};//{'a': 2, 'literal': 1, 'z': 2, 'op': 'addl'}
    instructions[3291] = {5'd2, 4'd0, 4'd2, 32'd9};//{'a': 2, 'b': 9, 'op': 'store'}
    instructions[3292] = {5'd0, 4'd8, 4'd0, 32'd65536};//{'literal': 65536, 'z': 8, 'op': 'literal'}
    instructions[3293] = {5'd0, 4'd9, 4'd0, 32'd0};//{'literal': 0, 'z': 9, 'op': 'literal'}
    instructions[3294] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3295] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3296] = {5'd2, 4'd0, 4'd3, 32'd9};//{'a': 3, 'comment': 'push', 'b': 9, 'op': 'store'}
    instructions[3297] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3298] = {5'd0, 4'd8, 4'd0, 32'd38};//{'literal': 38, 'z': 8, 'op': 'literal'}
    instructions[3299] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3300] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3301] = {5'd1, 4'd2, 4'd2, 32'd1};//{'a': 2, 'literal': 1, 'z': 2, 'op': 'addl'}
    instructions[3302] = {5'd5, 4'd9, 4'd2, 32'd0};//{'a': 2, 'z': 9, 'op': 'load'}
    instructions[3303] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3304] = {5'd5, 4'd11, 4'd3, 32'd0};//{'a': 3, 'z': 11, 'op': 'load'}
    instructions[3305] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3306] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[3307] = {5'd15, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'and'}
    instructions[3308] = {5'd15, 4'd9, 4'd9, 32'd11};//{'a': 9, 'z': 9, 'b': 11, 'op': 'and'}
    instructions[3309] = {5'd17, 4'd8, 4'd8, 32'd9};//{'a': 8, 'z': 8, 'b': 9, 'op': 'or'}
    instructions[3310] = {5'd6, 4'd0, 4'd8, 32'd3354};//{'a': 8, 'label': 3354, 'op': 'jmp_if_false'}
    instructions[3311] = {5'd0, 4'd8, 4'd0, 32'd65535};//{'literal': 65535, 'z': 8, 'op': 'literal'}
    instructions[3312] = {5'd0, 4'd9, 4'd0, 32'd0};//{'literal': 0, 'z': 9, 'op': 'literal'}
    instructions[3313] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3314] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3315] = {5'd2, 4'd0, 4'd3, 32'd9};//{'a': 3, 'comment': 'push', 'b': 9, 'op': 'store'}
    instructions[3316] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3317] = {5'd0, 4'd8, 4'd0, 32'd38};//{'literal': 38, 'z': 8, 'op': 'literal'}
    instructions[3318] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3319] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3320] = {5'd1, 4'd2, 4'd2, 32'd1};//{'a': 2, 'literal': 1, 'z': 2, 'op': 'addl'}
    instructions[3321] = {5'd5, 4'd9, 4'd2, 32'd0};//{'a': 2, 'z': 9, 'op': 'load'}
    instructions[3322] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3323] = {5'd5, 4'd11, 4'd3, 32'd0};//{'a': 3, 'z': 11, 'op': 'load'}
    instructions[3324] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3325] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[3326] = {5'd15, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'and'}
    instructions[3327] = {5'd15, 4'd9, 4'd9, 32'd11};//{'a': 9, 'z': 9, 'b': 11, 'op': 'and'}
    instructions[3328] = {5'd0, 4'd2, 4'd0, 32'd38};//{'literal': 38, 'z': 2, 'op': 'literal'}
    instructions[3329] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3330] = {5'd1, 4'd2, 4'd2, 32'd1};//{'a': 2, 'literal': 1, 'z': 2, 'op': 'addl'}
    instructions[3331] = {5'd2, 4'd0, 4'd2, 32'd9};//{'a': 2, 'b': 9, 'op': 'store'}
    instructions[3332] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[3333] = {5'd0, 4'd9, 4'd0, 32'd0};//{'literal': 0, 'z': 9, 'op': 'literal'}
    instructions[3334] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3335] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3336] = {5'd2, 4'd0, 4'd3, 32'd9};//{'a': 3, 'comment': 'push', 'b': 9, 'op': 'store'}
    instructions[3337] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3338] = {5'd0, 4'd8, 4'd0, 32'd38};//{'literal': 38, 'z': 8, 'op': 'literal'}
    instructions[3339] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3340] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3341] = {5'd1, 4'd2, 4'd2, 32'd1};//{'a': 2, 'literal': 1, 'z': 2, 'op': 'addl'}
    instructions[3342] = {5'd5, 4'd9, 4'd2, 32'd0};//{'a': 2, 'z': 9, 'op': 'load'}
    instructions[3343] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3344] = {5'd5, 4'd11, 4'd3, 32'd0};//{'a': 3, 'z': 11, 'op': 'load'}
    instructions[3345] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3346] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[3347] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[3348] = {5'd24, 4'd9, 4'd9, 32'd11};//{'a': 9, 'z': 9, 'b': 11, 'op': 'add_with_carry'}
    instructions[3349] = {5'd0, 4'd2, 4'd0, 32'd38};//{'literal': 38, 'z': 2, 'op': 'literal'}
    instructions[3350] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3351] = {5'd1, 4'd2, 4'd2, 32'd1};//{'a': 2, 'literal': 1, 'z': 2, 'op': 'addl'}
    instructions[3352] = {5'd2, 4'd0, 4'd2, 32'd9};//{'a': 2, 'b': 9, 'op': 'store'}
    instructions[3353] = {5'd8, 4'd0, 4'd0, 32'd3354};//{'label': 3354, 'op': 'goto'}
    instructions[3354] = {5'd1, 4'd3, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[3355] = {5'd1, 4'd4, 4'd7, 32'd0};//{'a': 7, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[3356] = {5'd12, 4'd0, 4'd6, 32'd0};//{'a': 6, 'op': 'return'}
    instructions[3357] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[3358] = {5'd0, 4'd8, 4'd0, 32'd38};//{'literal': 38, 'z': 8, 'op': 'literal'}
    instructions[3359] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3360] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3361] = {5'd1, 4'd2, 4'd2, 32'd1};//{'a': 2, 'literal': 1, 'z': 2, 'op': 'addl'}
    instructions[3362] = {5'd5, 4'd9, 4'd2, 32'd0};//{'a': 2, 'z': 9, 'op': 'load'}
    instructions[3363] = {5'd25, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'not'}
    instructions[3364] = {5'd25, 4'd9, 4'd9, 32'd0};//{'a': 9, 'z': 9, 'op': 'not'}
    instructions[3365] = {5'd0, 4'd2, 4'd0, 32'd43};//{'literal': 43, 'z': 2, 'op': 'literal'}
    instructions[3366] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3367] = {5'd1, 4'd3, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[3368] = {5'd1, 4'd4, 4'd7, 32'd0};//{'a': 7, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[3369] = {5'd12, 4'd0, 4'd6, 32'd0};//{'a': 6, 'op': 'return'}
    instructions[3370] = {5'd1, 4'd3, 4'd3, 32'd3};//{'a': 3, 'literal': 3, 'z': 3, 'op': 'addl'}
    instructions[3371] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[3372] = {5'd1, 4'd2, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3373] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3374] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[3375] = {5'd1, 4'd2, 4'd4, 32'd1};//{'a': 4, 'literal': 1, 'z': 2, 'op': 'addl'}
    instructions[3376] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3377] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[3378] = {5'd1, 4'd2, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 2, 'op': 'addl'}
    instructions[3379] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3380] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[3381] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3382] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[3383] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3384] = {5'd1, 4'd8, 4'd4, -32'd2};//{'a': 4, 'literal': -2, 'z': 8, 'op': 'addl'}
    instructions[3385] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3386] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3387] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3388] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3389] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[3390] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3391] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3392] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3393] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3394] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[3395] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[3396] = {5'd3, 4'd6, 4'd0, 32'd3762};//{'z': 6, 'label': 3762, 'op': 'call'}
    instructions[3397] = {5'd1, 4'd3, 4'd3, -32'd2};//{'a': 3, 'literal': -2, 'z': 3, 'op': 'addl'}
    instructions[3398] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3399] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[3400] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3401] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[3402] = {5'd0, 4'd2, 4'd0, 32'd2156};//{'literal': 2156, 'z': 2, 'op': 'literal'}
    instructions[3403] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3404] = {5'd1, 4'd2, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 2, 'op': 'addl'}
    instructions[3405] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3406] = {5'd0, 4'd8, 4'd0, 32'd17664};//{'literal': 17664, 'z': 8, 'op': 'literal'}
    instructions[3407] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3408] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3409] = {5'd1, 4'd8, 4'd4, -32'd5};//{'a': 4, 'literal': -5, 'z': 8, 'op': 'addl'}
    instructions[3410] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[3411] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3412] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3413] = {5'd0, 4'd8, 4'd0, 32'd7};//{'literal': 7, 'z': 8, 'op': 'literal'}
    instructions[3414] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3415] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[3416] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[3417] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3418] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3419] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[3420] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3421] = {5'd1, 4'd8, 4'd4, -32'd4};//{'a': 4, 'literal': -4, 'z': 8, 'op': 'addl'}
    instructions[3422] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3423] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3424] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3425] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3426] = {5'd1, 4'd8, 4'd4, -32'd5};//{'a': 4, 'literal': -5, 'z': 8, 'op': 'addl'}
    instructions[3427] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[3428] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3429] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3430] = {5'd0, 4'd8, 4'd0, 32'd8};//{'literal': 8, 'z': 8, 'op': 'literal'}
    instructions[3431] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3432] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[3433] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[3434] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3435] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3436] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[3437] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3438] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[3439] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3440] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3441] = {5'd1, 4'd8, 4'd4, -32'd5};//{'a': 4, 'literal': -5, 'z': 8, 'op': 'addl'}
    instructions[3442] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[3443] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3444] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3445] = {5'd0, 4'd8, 4'd0, 32'd9};//{'literal': 9, 'z': 8, 'op': 'literal'}
    instructions[3446] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3447] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[3448] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[3449] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3450] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3451] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[3452] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3453] = {5'd0, 4'd8, 4'd0, 32'd16384};//{'literal': 16384, 'z': 8, 'op': 'literal'}
    instructions[3454] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3455] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3456] = {5'd1, 4'd8, 4'd4, -32'd5};//{'a': 4, 'literal': -5, 'z': 8, 'op': 'addl'}
    instructions[3457] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[3458] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3459] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3460] = {5'd0, 4'd8, 4'd0, 32'd10};//{'literal': 10, 'z': 8, 'op': 'literal'}
    instructions[3461] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3462] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[3463] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[3464] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3465] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3466] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[3467] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3468] = {5'd1, 4'd8, 4'd4, -32'd3};//{'a': 4, 'literal': -3, 'z': 8, 'op': 'addl'}
    instructions[3469] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3470] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3471] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3472] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3473] = {5'd0, 4'd8, 4'd0, 32'd65280};//{'literal': 65280, 'z': 8, 'op': 'literal'}
    instructions[3474] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3475] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[3476] = {5'd17, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'or'}
    instructions[3477] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3478] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3479] = {5'd1, 4'd8, 4'd4, -32'd5};//{'a': 4, 'literal': -5, 'z': 8, 'op': 'addl'}
    instructions[3480] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[3481] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3482] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3483] = {5'd0, 4'd8, 4'd0, 32'd11};//{'literal': 11, 'z': 8, 'op': 'literal'}
    instructions[3484] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3485] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[3486] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[3487] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3488] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3489] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[3490] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3491] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[3492] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3493] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3494] = {5'd1, 4'd8, 4'd4, -32'd5};//{'a': 4, 'literal': -5, 'z': 8, 'op': 'addl'}
    instructions[3495] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[3496] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3497] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3498] = {5'd0, 4'd8, 4'd0, 32'd12};//{'literal': 12, 'z': 8, 'op': 'literal'}
    instructions[3499] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3500] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[3501] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[3502] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3503] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3504] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[3505] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3506] = {5'd0, 4'd8, 4'd0, 32'd49320};//{'literal': 49320, 'z': 8, 'op': 'literal'}
    instructions[3507] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3508] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3509] = {5'd1, 4'd8, 4'd4, -32'd5};//{'a': 4, 'literal': -5, 'z': 8, 'op': 'addl'}
    instructions[3510] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[3511] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3512] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3513] = {5'd0, 4'd8, 4'd0, 32'd13};//{'literal': 13, 'z': 8, 'op': 'literal'}
    instructions[3514] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3515] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[3516] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[3517] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3518] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3519] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[3520] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3521] = {5'd0, 4'd8, 4'd0, 32'd257};//{'literal': 257, 'z': 8, 'op': 'literal'}
    instructions[3522] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3523] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3524] = {5'd1, 4'd8, 4'd4, -32'd5};//{'a': 4, 'literal': -5, 'z': 8, 'op': 'addl'}
    instructions[3525] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[3526] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3527] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3528] = {5'd0, 4'd8, 4'd0, 32'd14};//{'literal': 14, 'z': 8, 'op': 'literal'}
    instructions[3529] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3530] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[3531] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[3532] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3533] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3534] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[3535] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3536] = {5'd1, 4'd8, 4'd4, -32'd2};//{'a': 4, 'literal': -2, 'z': 8, 'op': 'addl'}
    instructions[3537] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3538] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3539] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3540] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3541] = {5'd1, 4'd8, 4'd4, -32'd5};//{'a': 4, 'literal': -5, 'z': 8, 'op': 'addl'}
    instructions[3542] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[3543] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3544] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3545] = {5'd0, 4'd8, 4'd0, 32'd15};//{'literal': 15, 'z': 8, 'op': 'literal'}
    instructions[3546] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3547] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[3548] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[3549] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3550] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3551] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[3552] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3553] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[3554] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3555] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3556] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3557] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3558] = {5'd1, 4'd8, 4'd4, -32'd5};//{'a': 4, 'literal': -5, 'z': 8, 'op': 'addl'}
    instructions[3559] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[3560] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3561] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3562] = {5'd0, 4'd8, 4'd0, 32'd16};//{'literal': 16, 'z': 8, 'op': 'literal'}
    instructions[3563] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3564] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[3565] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[3566] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3567] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3568] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[3569] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3570] = {5'd0, 4'd8, 4'd0, 32'd14};//{'literal': 14, 'z': 8, 'op': 'literal'}
    instructions[3571] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3572] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3573] = {5'd1, 4'd8, 4'd4, -32'd4};//{'a': 4, 'literal': -4, 'z': 8, 'op': 'addl'}
    instructions[3574] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3575] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3576] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3577] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[3578] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[3579] = {5'd1, 4'd2, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3580] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3581] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[3582] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3583] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[3584] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3585] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[3586] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[3587] = {5'd3, 4'd6, 4'd0, 32'd3258};//{'z': 6, 'label': 3258, 'op': 'call'}
    instructions[3588] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[3589] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3590] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[3591] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3592] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[3593] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[3594] = {5'd0, 4'd8, 4'd0, 32'd7};//{'literal': 7, 'z': 8, 'op': 'literal'}
    instructions[3595] = {5'd1, 4'd2, 4'd4, 32'd1};//{'a': 4, 'literal': 1, 'z': 2, 'op': 'addl'}
    instructions[3596] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3597] = {5'd1, 4'd8, 4'd4, 32'd1};//{'a': 4, 'literal': 1, 'z': 8, 'op': 'addl'}
    instructions[3598] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3599] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3600] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3601] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3602] = {5'd0, 4'd8, 4'd0, 32'd16};//{'literal': 16, 'z': 8, 'op': 'literal'}
    instructions[3603] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3604] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[3605] = {5'd19, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'unsigned_greater_equal'}
    instructions[3606] = {5'd6, 4'd0, 4'd8, 32'd3653};//{'a': 8, 'label': 3653, 'op': 'jmp_if_false'}
    instructions[3607] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[3608] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3609] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[3610] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3611] = {5'd1, 4'd8, 4'd4, -32'd5};//{'a': 4, 'literal': -5, 'z': 8, 'op': 'addl'}
    instructions[3612] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[3613] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3614] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3615] = {5'd1, 4'd8, 4'd4, 32'd1};//{'a': 4, 'literal': 1, 'z': 8, 'op': 'addl'}
    instructions[3616] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3617] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3618] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3619] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[3620] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[3621] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3622] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3623] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3624] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3625] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[3626] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[3627] = {5'd3, 4'd6, 4'd0, 32'd3268};//{'z': 6, 'label': 3268, 'op': 'call'}
    instructions[3628] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3629] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3630] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[3631] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3632] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[3633] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[3634] = {5'd1, 4'd8, 4'd4, 32'd1};//{'a': 4, 'literal': 1, 'z': 8, 'op': 'addl'}
    instructions[3635] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3636] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3637] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3638] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3639] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[3640] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3641] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3642] = {5'd1, 4'd8, 4'd4, 32'd1};//{'a': 4, 'literal': 1, 'z': 8, 'op': 'addl'}
    instructions[3643] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3644] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3645] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3646] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[3647] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[3648] = {5'd1, 4'd2, 4'd4, 32'd1};//{'a': 4, 'literal': 1, 'z': 2, 'op': 'addl'}
    instructions[3649] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3650] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3651] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[3652] = {5'd8, 4'd0, 4'd0, 32'd3597};//{'label': 3597, 'op': 'goto'}
    instructions[3653] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[3654] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3655] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[3656] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3657] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[3658] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[3659] = {5'd3, 4'd6, 4'd0, 32'd3357};//{'z': 6, 'label': 3357, 'op': 'call'}
    instructions[3660] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[3661] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3662] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[3663] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3664] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[3665] = {5'd0, 4'd2, 4'd0, 32'd43};//{'literal': 43, 'z': 2, 'op': 'literal'}
    instructions[3666] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3667] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3668] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3669] = {5'd1, 4'd8, 4'd4, -32'd5};//{'a': 4, 'literal': -5, 'z': 8, 'op': 'addl'}
    instructions[3670] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[3671] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3672] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3673] = {5'd0, 4'd8, 4'd0, 32'd12};//{'literal': 12, 'z': 8, 'op': 'literal'}
    instructions[3674] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3675] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[3676] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[3677] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3678] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3679] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[3680] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3681] = {5'd1, 4'd8, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 8, 'op': 'addl'}
    instructions[3682] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3683] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3684] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3685] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3686] = {5'd0, 4'd8, 4'd0, 32'd64};//{'literal': 64, 'z': 8, 'op': 'literal'}
    instructions[3687] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3688] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[3689] = {5'd20, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'unsigned_greater'}
    instructions[3690] = {5'd6, 4'd0, 4'd8, 32'd3695};//{'a': 8, 'label': 3695, 'op': 'jmp_if_false'}
    instructions[3691] = {5'd0, 4'd8, 4'd0, 32'd64};//{'literal': 64, 'z': 8, 'op': 'literal'}
    instructions[3692] = {5'd1, 4'd2, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3693] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3694] = {5'd8, 4'd0, 4'd0, 32'd3695};//{'label': 3695, 'op': 'goto'}
    instructions[3695] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[3696] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3697] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[3698] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3699] = {5'd1, 4'd8, 4'd4, -32'd5};//{'a': 4, 'literal': -5, 'z': 8, 'op': 'addl'}
    instructions[3700] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[3701] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3702] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3703] = {5'd1, 4'd8, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 8, 'op': 'addl'}
    instructions[3704] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3705] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3706] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3707] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3708] = {5'd0, 4'd8, 4'd0, 32'd2705};//{'literal': 2705, 'z': 8, 'op': 'literal'}
    instructions[3709] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3710] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3711] = {5'd1, 4'd8, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 8, 'op': 'addl'}
    instructions[3712] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3713] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3714] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3715] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[3716] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[3717] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3718] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3719] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3720] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3721] = {5'd0, 4'd8, 4'd0, 32'd2728};//{'literal': 2728, 'z': 8, 'op': 'literal'}
    instructions[3722] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3723] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3724] = {5'd1, 4'd8, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 8, 'op': 'addl'}
    instructions[3725] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3726] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3727] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3728] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[3729] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[3730] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3731] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3732] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3733] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3734] = {5'd0, 4'd8, 4'd0, 32'd1093};//{'literal': 1093, 'z': 8, 'op': 'literal'}
    instructions[3735] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3736] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3737] = {5'd1, 4'd8, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 8, 'op': 'addl'}
    instructions[3738] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3739] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3740] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3741] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[3742] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[3743] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3744] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3745] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3746] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3747] = {5'd0, 4'd8, 4'd0, 32'd2048};//{'literal': 2048, 'z': 8, 'op': 'literal'}
    instructions[3748] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3749] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3750] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[3751] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[3752] = {5'd3, 4'd6, 4'd0, 32'd3026};//{'z': 6, 'label': 3026, 'op': 'call'}
    instructions[3753] = {5'd1, 4'd3, 4'd3, -32'd6};//{'a': 3, 'literal': -6, 'z': 3, 'op': 'addl'}
    instructions[3754] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3755] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[3756] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3757] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[3758] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[3759] = {5'd1, 4'd3, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[3760] = {5'd1, 4'd4, 4'd7, 32'd0};//{'a': 7, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[3761] = {5'd12, 4'd0, 4'd6, 32'd0};//{'a': 6, 'op': 'return'}
    instructions[3762] = {5'd1, 4'd3, 4'd3, 32'd19};//{'a': 3, 'literal': 19, 'z': 3, 'op': 'addl'}
    instructions[3763] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[3764] = {5'd1, 4'd2, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3765] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3766] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[3767] = {5'd1, 4'd2, 4'd4, 32'd1};//{'a': 4, 'literal': 1, 'z': 2, 'op': 'addl'}
    instructions[3768] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3769] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[3770] = {5'd1, 4'd2, 4'd4, 32'd18};//{'a': 4, 'literal': 18, 'z': 2, 'op': 'addl'}
    instructions[3771] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3772] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[3773] = {5'd1, 4'd2, 4'd4, 32'd18};//{'a': 4, 'literal': 18, 'z': 2, 'op': 'addl'}
    instructions[3774] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3775] = {5'd1, 4'd8, 4'd4, 32'd18};//{'a': 4, 'literal': 18, 'z': 8, 'op': 'addl'}
    instructions[3776] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3777] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3778] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3779] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3780] = {5'd0, 4'd8, 4'd0, 32'd16};//{'literal': 16, 'z': 8, 'op': 'literal'}
    instructions[3781] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3782] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[3783] = {5'd20, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'unsigned_greater'}
    instructions[3784] = {5'd6, 4'd0, 4'd8, 32'd3853};//{'a': 8, 'label': 3853, 'op': 'jmp_if_false'}
    instructions[3785] = {5'd1, 4'd8, 4'd4, -32'd2};//{'a': 4, 'literal': -2, 'z': 8, 'op': 'addl'}
    instructions[3786] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3787] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3788] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3789] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3790] = {5'd0, 4'd8, 4'd0, 32'd17};//{'literal': 17, 'z': 8, 'op': 'literal'}
    instructions[3791] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3792] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3793] = {5'd1, 4'd8, 4'd4, 32'd18};//{'a': 4, 'literal': 18, 'z': 8, 'op': 'addl'}
    instructions[3794] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3795] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3796] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3797] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[3798] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[3799] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3800] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3801] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3802] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[3803] = {5'd7, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'equal'}
    instructions[3804] = {5'd6, 4'd0, 4'd8, 32'd3824};//{'a': 8, 'label': 3824, 'op': 'jmp_if_false'}
    instructions[3805] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[3806] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3807] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3808] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3809] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3810] = {5'd0, 4'd8, 4'd0, 32'd2157};//{'literal': 2157, 'z': 8, 'op': 'literal'}
    instructions[3811] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3812] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3813] = {5'd1, 4'd8, 4'd4, 32'd18};//{'a': 4, 'literal': 18, 'z': 8, 'op': 'addl'}
    instructions[3814] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3815] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3816] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3817] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[3818] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[3819] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3820] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3821] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3822] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[3823] = {5'd7, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'equal'}
    instructions[3824] = {5'd6, 4'd0, 4'd8, 32'd3834};//{'a': 8, 'label': 3834, 'op': 'jmp_if_false'}
    instructions[3825] = {5'd1, 4'd8, 4'd4, 32'd18};//{'a': 4, 'literal': 18, 'z': 8, 'op': 'addl'}
    instructions[3826] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3827] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3828] = {5'd0, 4'd2, 4'd0, 32'd2156};//{'literal': 2156, 'z': 2, 'op': 'literal'}
    instructions[3829] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3830] = {5'd1, 4'd3, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[3831] = {5'd1, 4'd4, 4'd7, 32'd0};//{'a': 7, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[3832] = {5'd12, 4'd0, 4'd6, 32'd0};//{'a': 6, 'op': 'return'}
    instructions[3833] = {5'd8, 4'd0, 4'd0, 32'd3834};//{'label': 3834, 'op': 'goto'}
    instructions[3834] = {5'd1, 4'd8, 4'd4, 32'd18};//{'a': 4, 'literal': 18, 'z': 8, 'op': 'addl'}
    instructions[3835] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3836] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3837] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3838] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3839] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[3840] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3841] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3842] = {5'd1, 4'd8, 4'd4, 32'd18};//{'a': 4, 'literal': 18, 'z': 8, 'op': 'addl'}
    instructions[3843] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3844] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3845] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3846] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[3847] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[3848] = {5'd1, 4'd2, 4'd4, 32'd18};//{'a': 4, 'literal': 18, 'z': 2, 'op': 'addl'}
    instructions[3849] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3850] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3851] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[3852] = {5'd8, 4'd0, 4'd0, 32'd3775};//{'label': 3775, 'op': 'goto'}
    instructions[3853] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[3854] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3855] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3856] = {5'd0, 4'd8, 4'd0, 32'd2173};//{'literal': 2173, 'z': 8, 'op': 'literal'}
    instructions[3857] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3858] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3859] = {5'd0, 4'd8, 4'd0, 32'd7};//{'literal': 7, 'z': 8, 'op': 'literal'}
    instructions[3860] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3861] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[3862] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[3863] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3864] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3865] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[3866] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3867] = {5'd0, 4'd8, 4'd0, 32'd2048};//{'literal': 2048, 'z': 8, 'op': 'literal'}
    instructions[3868] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3869] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3870] = {5'd0, 4'd8, 4'd0, 32'd2173};//{'literal': 2173, 'z': 8, 'op': 'literal'}
    instructions[3871] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3872] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3873] = {5'd0, 4'd8, 4'd0, 32'd8};//{'literal': 8, 'z': 8, 'op': 'literal'}
    instructions[3874] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3875] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[3876] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[3877] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3878] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3879] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[3880] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3881] = {5'd0, 4'd8, 4'd0, 32'd1540};//{'literal': 1540, 'z': 8, 'op': 'literal'}
    instructions[3882] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3883] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3884] = {5'd0, 4'd8, 4'd0, 32'd2173};//{'literal': 2173, 'z': 8, 'op': 'literal'}
    instructions[3885] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3886] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3887] = {5'd0, 4'd8, 4'd0, 32'd9};//{'literal': 9, 'z': 8, 'op': 'literal'}
    instructions[3888] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3889] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[3890] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[3891] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3892] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3893] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[3894] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3895] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[3896] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3897] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3898] = {5'd0, 4'd8, 4'd0, 32'd2173};//{'literal': 2173, 'z': 8, 'op': 'literal'}
    instructions[3899] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3900] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3901] = {5'd0, 4'd8, 4'd0, 32'd10};//{'literal': 10, 'z': 8, 'op': 'literal'}
    instructions[3902] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3903] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[3904] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[3905] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3906] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3907] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[3908] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3909] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[3910] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3911] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3912] = {5'd0, 4'd8, 4'd0, 32'd2173};//{'literal': 2173, 'z': 8, 'op': 'literal'}
    instructions[3913] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3914] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3915] = {5'd0, 4'd8, 4'd0, 32'd11};//{'literal': 11, 'z': 8, 'op': 'literal'}
    instructions[3916] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3917] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[3918] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[3919] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3920] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3921] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[3922] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3923] = {5'd0, 4'd8, 4'd0, 32'd515};//{'literal': 515, 'z': 8, 'op': 'literal'}
    instructions[3924] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3925] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3926] = {5'd0, 4'd8, 4'd0, 32'd2173};//{'literal': 2173, 'z': 8, 'op': 'literal'}
    instructions[3927] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3928] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3929] = {5'd0, 4'd8, 4'd0, 32'd12};//{'literal': 12, 'z': 8, 'op': 'literal'}
    instructions[3930] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3931] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[3932] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[3933] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3934] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3935] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[3936] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3937] = {5'd0, 4'd8, 4'd0, 32'd1029};//{'literal': 1029, 'z': 8, 'op': 'literal'}
    instructions[3938] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3939] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3940] = {5'd0, 4'd8, 4'd0, 32'd2173};//{'literal': 2173, 'z': 8, 'op': 'literal'}
    instructions[3941] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3942] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3943] = {5'd0, 4'd8, 4'd0, 32'd13};//{'literal': 13, 'z': 8, 'op': 'literal'}
    instructions[3944] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3945] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[3946] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[3947] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3948] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3949] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[3950] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3951] = {5'd0, 4'd8, 4'd0, 32'd49320};//{'literal': 49320, 'z': 8, 'op': 'literal'}
    instructions[3952] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3953] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3954] = {5'd0, 4'd8, 4'd0, 32'd2173};//{'literal': 2173, 'z': 8, 'op': 'literal'}
    instructions[3955] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3956] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3957] = {5'd0, 4'd8, 4'd0, 32'd14};//{'literal': 14, 'z': 8, 'op': 'literal'}
    instructions[3958] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3959] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[3960] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[3961] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3962] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3963] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[3964] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3965] = {5'd0, 4'd8, 4'd0, 32'd257};//{'literal': 257, 'z': 8, 'op': 'literal'}
    instructions[3966] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3967] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3968] = {5'd0, 4'd8, 4'd0, 32'd2173};//{'literal': 2173, 'z': 8, 'op': 'literal'}
    instructions[3969] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3970] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3971] = {5'd0, 4'd8, 4'd0, 32'd15};//{'literal': 15, 'z': 8, 'op': 'literal'}
    instructions[3972] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3973] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[3974] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[3975] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3976] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3977] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[3978] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3979] = {5'd1, 4'd8, 4'd4, -32'd2};//{'a': 4, 'literal': -2, 'z': 8, 'op': 'addl'}
    instructions[3980] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3981] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3982] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3983] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3984] = {5'd0, 4'd8, 4'd0, 32'd2173};//{'literal': 2173, 'z': 8, 'op': 'literal'}
    instructions[3985] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3986] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[3987] = {5'd0, 4'd8, 4'd0, 32'd19};//{'literal': 19, 'z': 8, 'op': 'literal'}
    instructions[3988] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3989] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[3990] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[3991] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3992] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[3993] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[3994] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[3995] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[3996] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[3997] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[3998] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[3999] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4000] = {5'd0, 4'd8, 4'd0, 32'd2173};//{'literal': 2173, 'z': 8, 'op': 'literal'}
    instructions[4001] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4002] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4003] = {5'd0, 4'd8, 4'd0, 32'd20};//{'literal': 20, 'z': 8, 'op': 'literal'}
    instructions[4004] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4005] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[4006] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[4007] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4008] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4009] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[4010] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[4011] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[4012] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4013] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[4014] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4015] = {5'd0, 4'd8, 4'd0, 32'd2173};//{'literal': 2173, 'z': 8, 'op': 'literal'}
    instructions[4016] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4017] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4018] = {5'd0, 4'd8, 4'd0, 32'd64};//{'literal': 64, 'z': 8, 'op': 'literal'}
    instructions[4019] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4020] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4021] = {5'd0, 4'd8, 4'd0, 32'd65535};//{'literal': 65535, 'z': 8, 'op': 'literal'}
    instructions[4022] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4023] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4024] = {5'd0, 4'd8, 4'd0, 32'd65535};//{'literal': 65535, 'z': 8, 'op': 'literal'}
    instructions[4025] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4026] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4027] = {5'd0, 4'd8, 4'd0, 32'd65535};//{'literal': 65535, 'z': 8, 'op': 'literal'}
    instructions[4028] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4029] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4030] = {5'd0, 4'd8, 4'd0, 32'd2054};//{'literal': 2054, 'z': 8, 'op': 'literal'}
    instructions[4031] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4032] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4033] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[4034] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[4035] = {5'd3, 4'd6, 4'd0, 32'd3026};//{'z': 6, 'label': 3026, 'op': 'call'}
    instructions[4036] = {5'd1, 4'd3, 4'd3, -32'd6};//{'a': 3, 'literal': -6, 'z': 3, 'op': 'addl'}
    instructions[4037] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4038] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[4039] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4040] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[4041] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[4042] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[4043] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4044] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[4045] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4046] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[4047] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[4048] = {5'd3, 4'd6, 4'd0, 32'd3016};//{'z': 6, 'label': 3016, 'op': 'call'}
    instructions[4049] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[4050] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4051] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[4052] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4053] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[4054] = {5'd0, 4'd2, 4'd0, 32'd1081};//{'literal': 1081, 'z': 2, 'op': 'literal'}
    instructions[4055] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4056] = {5'd1, 4'd2, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4057] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[4058] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[4059] = {5'd1, 4'd2, 4'd4, 32'd18};//{'a': 4, 'literal': 18, 'z': 2, 'op': 'addl'}
    instructions[4060] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[4061] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[4062] = {5'd1, 4'd2, 4'd4, 32'd1};//{'a': 4, 'literal': 1, 'z': 2, 'op': 'addl'}
    instructions[4063] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[4064] = {5'd1, 4'd8, 4'd4, 32'd1};//{'a': 4, 'literal': 1, 'z': 8, 'op': 'addl'}
    instructions[4065] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4066] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4067] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4068] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4069] = {5'd1, 4'd8, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 8, 'op': 'addl'}
    instructions[4070] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4071] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4072] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4073] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[4074] = {5'd20, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'unsigned_greater'}
    instructions[4075] = {5'd6, 4'd0, 4'd8, 32'd4160};//{'a': 8, 'label': 4160, 'op': 'jmp_if_false'}
    instructions[4076] = {5'd1, 4'd8, 4'd4, 32'd18};//{'a': 4, 'literal': 18, 'z': 8, 'op': 'addl'}
    instructions[4077] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4078] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4079] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4080] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4081] = {5'd0, 4'd8, 4'd0, 32'd16};//{'literal': 16, 'z': 8, 'op': 'literal'}
    instructions[4082] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4083] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[4084] = {5'd20, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'unsigned_greater'}
    instructions[4085] = {5'd6, 4'd0, 4'd8, 32'd4116};//{'a': 8, 'label': 4116, 'op': 'jmp_if_false'}
    instructions[4086] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[4087] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4088] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[4089] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4090] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[4091] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[4092] = {5'd3, 4'd6, 4'd0, 32'd3016};//{'z': 6, 'label': 3016, 'op': 'call'}
    instructions[4093] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[4094] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4095] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[4096] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4097] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[4098] = {5'd0, 4'd2, 4'd0, 32'd1081};//{'literal': 1081, 'z': 2, 'op': 'literal'}
    instructions[4099] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4100] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4101] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4102] = {5'd1, 4'd8, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 8, 'op': 'addl'}
    instructions[4103] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4104] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4105] = {5'd1, 4'd8, 4'd4, 32'd18};//{'a': 4, 'literal': 18, 'z': 8, 'op': 'addl'}
    instructions[4106] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4107] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4108] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4109] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[4110] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[4111] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4112] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4113] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[4114] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[4115] = {5'd8, 4'd0, 4'd0, 32'd4130};//{'label': 4130, 'op': 'goto'}
    instructions[4116] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[4117] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4118] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[4119] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4120] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[4121] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[4122] = {5'd3, 4'd6, 4'd0, 32'd3016};//{'z': 6, 'label': 3016, 'op': 'call'}
    instructions[4123] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[4124] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4125] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[4126] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4127] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[4128] = {5'd0, 4'd2, 4'd0, 32'd1081};//{'literal': 1081, 'z': 2, 'op': 'literal'}
    instructions[4129] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4130] = {5'd1, 4'd8, 4'd4, 32'd18};//{'a': 4, 'literal': 18, 'z': 8, 'op': 'addl'}
    instructions[4131] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4132] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4133] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4134] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4135] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[4136] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4137] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4138] = {5'd1, 4'd8, 4'd4, 32'd18};//{'a': 4, 'literal': 18, 'z': 8, 'op': 'addl'}
    instructions[4139] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4140] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4141] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4142] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[4143] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[4144] = {5'd1, 4'd2, 4'd4, 32'd18};//{'a': 4, 'literal': 18, 'z': 2, 'op': 'addl'}
    instructions[4145] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[4146] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4147] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[4148] = {5'd0, 4'd8, 4'd0, 32'd2};//{'literal': 2, 'z': 8, 'op': 'literal'}
    instructions[4149] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4150] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4151] = {5'd1, 4'd8, 4'd4, 32'd1};//{'a': 4, 'literal': 1, 'z': 8, 'op': 'addl'}
    instructions[4152] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4153] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4154] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4155] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[4156] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[4157] = {5'd1, 4'd2, 4'd4, 32'd1};//{'a': 4, 'literal': 1, 'z': 2, 'op': 'addl'}
    instructions[4158] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[4159] = {5'd8, 4'd0, 4'd0, 32'd4064};//{'label': 4064, 'op': 'goto'}
    instructions[4160] = {5'd0, 4'd8, 4'd0, 32'd2054};//{'literal': 2054, 'z': 8, 'op': 'literal'}
    instructions[4161] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4162] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4163] = {5'd1, 4'd8, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 8, 'op': 'addl'}
    instructions[4164] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4165] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4166] = {5'd0, 4'd8, 4'd0, 32'd6};//{'literal': 6, 'z': 8, 'op': 'literal'}
    instructions[4167] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4168] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[4169] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[4170] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4171] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4172] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4173] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[4174] = {5'd7, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'equal'}
    instructions[4175] = {5'd6, 4'd0, 4'd8, 32'd4191};//{'a': 8, 'label': 4191, 'op': 'jmp_if_false'}
    instructions[4176] = {5'd0, 4'd8, 4'd0, 32'd2};//{'literal': 2, 'z': 8, 'op': 'literal'}
    instructions[4177] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4178] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4179] = {5'd1, 4'd8, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 8, 'op': 'addl'}
    instructions[4180] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4181] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4182] = {5'd0, 4'd8, 4'd0, 32'd10};//{'literal': 10, 'z': 8, 'op': 'literal'}
    instructions[4183] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4184] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[4185] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[4186] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4187] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4188] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4189] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[4190] = {5'd7, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'equal'}
    instructions[4191] = {5'd6, 4'd0, 4'd8, 32'd4383};//{'a': 8, 'label': 4383, 'op': 'jmp_if_false'}
    instructions[4192] = {5'd1, 4'd8, 4'd4, -32'd2};//{'a': 4, 'literal': -2, 'z': 8, 'op': 'addl'}
    instructions[4193] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4194] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4195] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4196] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4197] = {5'd1, 4'd8, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 8, 'op': 'addl'}
    instructions[4198] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4199] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4200] = {5'd0, 4'd8, 4'd0, 32'd14};//{'literal': 14, 'z': 8, 'op': 'literal'}
    instructions[4201] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4202] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[4203] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[4204] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4205] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4206] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4207] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[4208] = {5'd7, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'equal'}
    instructions[4209] = {5'd6, 4'd0, 4'd8, 32'd4227};//{'a': 8, 'label': 4227, 'op': 'jmp_if_false'}
    instructions[4210] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[4211] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4212] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4213] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4214] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4215] = {5'd1, 4'd8, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 8, 'op': 'addl'}
    instructions[4216] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4217] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4218] = {5'd0, 4'd8, 4'd0, 32'd15};//{'literal': 15, 'z': 8, 'op': 'literal'}
    instructions[4219] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4220] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[4221] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[4222] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4223] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4224] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4225] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[4226] = {5'd7, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'equal'}
    instructions[4227] = {5'd6, 4'd0, 4'd8, 32'd4382};//{'a': 8, 'label': 4382, 'op': 'jmp_if_false'}
    instructions[4228] = {5'd1, 4'd8, 4'd4, -32'd2};//{'a': 4, 'literal': -2, 'z': 8, 'op': 'addl'}
    instructions[4229] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4230] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4231] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4232] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4233] = {5'd0, 4'd8, 4'd0, 32'd17};//{'literal': 17, 'z': 8, 'op': 'literal'}
    instructions[4234] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4235] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4236] = {5'd0, 4'd8, 4'd0, 32'd37};//{'literal': 37, 'z': 8, 'op': 'literal'}
    instructions[4237] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4238] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4239] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4240] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[4241] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[4242] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4243] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4244] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[4245] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[4246] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[4247] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4248] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4249] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4250] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4251] = {5'd0, 4'd8, 4'd0, 32'd2157};//{'literal': 2157, 'z': 8, 'op': 'literal'}
    instructions[4252] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4253] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4254] = {5'd0, 4'd8, 4'd0, 32'd37};//{'literal': 37, 'z': 8, 'op': 'literal'}
    instructions[4255] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4256] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4257] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4258] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[4259] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[4260] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4261] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4262] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[4263] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[4264] = {5'd1, 4'd8, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 8, 'op': 'addl'}
    instructions[4265] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4266] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4267] = {5'd0, 4'd8, 4'd0, 32'd11};//{'literal': 11, 'z': 8, 'op': 'literal'}
    instructions[4268] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4269] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[4270] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[4271] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4272] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4273] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4274] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4275] = {5'd0, 4'd8, 4'd0, 32'd2705};//{'literal': 2705, 'z': 8, 'op': 'literal'}
    instructions[4276] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4277] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4278] = {5'd0, 4'd8, 4'd0, 32'd37};//{'literal': 37, 'z': 8, 'op': 'literal'}
    instructions[4279] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4280] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4281] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4282] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[4283] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[4284] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4285] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4286] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[4287] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[4288] = {5'd1, 4'd8, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 8, 'op': 'addl'}
    instructions[4289] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4290] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4291] = {5'd0, 4'd8, 4'd0, 32'd12};//{'literal': 12, 'z': 8, 'op': 'literal'}
    instructions[4292] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4293] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[4294] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[4295] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4296] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4297] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4298] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4299] = {5'd0, 4'd8, 4'd0, 32'd2728};//{'literal': 2728, 'z': 8, 'op': 'literal'}
    instructions[4300] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4301] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4302] = {5'd0, 4'd8, 4'd0, 32'd37};//{'literal': 37, 'z': 8, 'op': 'literal'}
    instructions[4303] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4304] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4305] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4306] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[4307] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[4308] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4309] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4310] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[4311] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[4312] = {5'd1, 4'd8, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 8, 'op': 'addl'}
    instructions[4313] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4314] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4315] = {5'd0, 4'd8, 4'd0, 32'd13};//{'literal': 13, 'z': 8, 'op': 'literal'}
    instructions[4316] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4317] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[4318] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[4319] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4320] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4321] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4322] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4323] = {5'd0, 4'd8, 4'd0, 32'd1093};//{'literal': 1093, 'z': 8, 'op': 'literal'}
    instructions[4324] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4325] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4326] = {5'd0, 4'd8, 4'd0, 32'd37};//{'literal': 37, 'z': 8, 'op': 'literal'}
    instructions[4327] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4328] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4329] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4330] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[4331] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[4332] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4333] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4334] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[4335] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[4336] = {5'd0, 4'd8, 4'd0, 32'd37};//{'literal': 37, 'z': 8, 'op': 'literal'}
    instructions[4337] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4338] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4339] = {5'd1, 4'd2, 4'd4, 32'd18};//{'a': 4, 'literal': 18, 'z': 2, 'op': 'addl'}
    instructions[4340] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[4341] = {5'd0, 4'd8, 4'd0, 32'd37};//{'literal': 37, 'z': 8, 'op': 'literal'}
    instructions[4342] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4343] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4344] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4345] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4346] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[4347] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4348] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4349] = {5'd0, 4'd8, 4'd0, 32'd37};//{'literal': 37, 'z': 8, 'op': 'literal'}
    instructions[4350] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4351] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4352] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4353] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[4354] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[4355] = {5'd0, 4'd2, 4'd0, 32'd37};//{'literal': 37, 'z': 2, 'op': 'literal'}
    instructions[4356] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[4357] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4358] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[4359] = {5'd0, 4'd8, 4'd0, 32'd16};//{'literal': 16, 'z': 8, 'op': 'literal'}
    instructions[4360] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4361] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4362] = {5'd0, 4'd8, 4'd0, 32'd37};//{'literal': 37, 'z': 8, 'op': 'literal'}
    instructions[4363] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4364] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4365] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4366] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[4367] = {5'd7, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'equal'}
    instructions[4368] = {5'd6, 4'd0, 4'd8, 32'd4373};//{'a': 8, 'label': 4373, 'op': 'jmp_if_false'}
    instructions[4369] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[4370] = {5'd0, 4'd2, 4'd0, 32'd37};//{'literal': 37, 'z': 2, 'op': 'literal'}
    instructions[4371] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[4372] = {5'd8, 4'd0, 4'd0, 32'd4373};//{'label': 4373, 'op': 'goto'}
    instructions[4373] = {5'd1, 4'd8, 4'd4, 32'd18};//{'a': 4, 'literal': 18, 'z': 8, 'op': 'addl'}
    instructions[4374] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4375] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4376] = {5'd0, 4'd2, 4'd0, 32'd2156};//{'literal': 2156, 'z': 2, 'op': 'literal'}
    instructions[4377] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[4378] = {5'd1, 4'd3, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[4379] = {5'd1, 4'd4, 4'd7, 32'd0};//{'a': 7, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[4380] = {5'd12, 4'd0, 4'd6, 32'd0};//{'a': 6, 'op': 'return'}
    instructions[4381] = {5'd8, 4'd0, 4'd0, 32'd4382};//{'label': 4382, 'op': 'goto'}
    instructions[4382] = {5'd8, 4'd0, 4'd0, 32'd4383};//{'label': 4383, 'op': 'goto'}
    instructions[4383] = {5'd8, 4'd0, 4'd0, 32'd4042};//{'label': 4042, 'op': 'goto'}
    instructions[4384] = {5'd1, 4'd3, 4'd3, 32'd4};//{'a': 3, 'literal': 4, 'z': 3, 'op': 'addl'}
    instructions[4385] = {5'd0, 4'd8, 4'd0, 32'd17};//{'literal': 17, 'z': 8, 'op': 'literal'}
    instructions[4386] = {5'd1, 4'd2, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4387] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[4388] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[4389] = {5'd1, 4'd2, 4'd4, 32'd1};//{'a': 4, 'literal': 1, 'z': 2, 'op': 'addl'}
    instructions[4390] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[4391] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[4392] = {5'd1, 4'd2, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 2, 'op': 'addl'}
    instructions[4393] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[4394] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[4395] = {5'd1, 4'd2, 4'd4, 32'd3};//{'a': 4, 'literal': 3, 'z': 2, 'op': 'addl'}
    instructions[4396] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[4397] = {5'd0, 4'd8, 4'd0, 32'd1091};//{'literal': 1091, 'z': 8, 'op': 'literal'}
    instructions[4398] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4399] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4400] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4401] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4402] = {5'd1, 4'd8, 4'd4, -32'd2};//{'a': 4, 'literal': -2, 'z': 8, 'op': 'addl'}
    instructions[4403] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[4404] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4405] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4406] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[4407] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4408] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4409] = {5'd1, 4'd8, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 8, 'op': 'addl'}
    instructions[4410] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4411] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4412] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4413] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[4414] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[4415] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4416] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[4417] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[4418] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4419] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4420] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[4421] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[4422] = {5'd0, 4'd8, 4'd0, 32'd1078};//{'literal': 1078, 'z': 8, 'op': 'literal'}
    instructions[4423] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4424] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4425] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4426] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4427] = {5'd1, 4'd8, 4'd4, -32'd2};//{'a': 4, 'literal': -2, 'z': 8, 'op': 'addl'}
    instructions[4428] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[4429] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4430] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4431] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[4432] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4433] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4434] = {5'd1, 4'd8, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 8, 'op': 'addl'}
    instructions[4435] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4436] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4437] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4438] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[4439] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[4440] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4441] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[4442] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[4443] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4444] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4445] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[4446] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[4447] = {5'd0, 4'd8, 4'd0, 32'd16};//{'literal': 16, 'z': 8, 'op': 'literal'}
    instructions[4448] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4449] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4450] = {5'd0, 4'd8, 4'd0, 32'd2703};//{'literal': 2703, 'z': 8, 'op': 'literal'}
    instructions[4451] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4452] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4453] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4454] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[4455] = {5'd14, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'unsigned_shift_right'}
    instructions[4456] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4457] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4458] = {5'd1, 4'd8, 4'd4, -32'd2};//{'a': 4, 'literal': -2, 'z': 8, 'op': 'addl'}
    instructions[4459] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[4460] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4461] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4462] = {5'd0, 4'd8, 4'd0, 32'd2};//{'literal': 2, 'z': 8, 'op': 'literal'}
    instructions[4463] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4464] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4465] = {5'd1, 4'd8, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 8, 'op': 'addl'}
    instructions[4466] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4467] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4468] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4469] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[4470] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[4471] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4472] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[4473] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[4474] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4475] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4476] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[4477] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[4478] = {5'd0, 4'd8, 4'd0, 32'd65535};//{'literal': 65535, 'z': 8, 'op': 'literal'}
    instructions[4479] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4480] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4481] = {5'd0, 4'd8, 4'd0, 32'd2703};//{'literal': 2703, 'z': 8, 'op': 'literal'}
    instructions[4482] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4483] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4484] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4485] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[4486] = {5'd15, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'and'}
    instructions[4487] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4488] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4489] = {5'd1, 4'd8, 4'd4, -32'd2};//{'a': 4, 'literal': -2, 'z': 8, 'op': 'addl'}
    instructions[4490] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[4491] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4492] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4493] = {5'd0, 4'd8, 4'd0, 32'd3};//{'literal': 3, 'z': 8, 'op': 'literal'}
    instructions[4494] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4495] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4496] = {5'd1, 4'd8, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 8, 'op': 'addl'}
    instructions[4497] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4498] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4499] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4500] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[4501] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[4502] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4503] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[4504] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[4505] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4506] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4507] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[4508] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[4509] = {5'd0, 4'd8, 4'd0, 32'd16};//{'literal': 16, 'z': 8, 'op': 'literal'}
    instructions[4510] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4511] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4512] = {5'd0, 4'd8, 4'd0, 32'd46};//{'literal': 46, 'z': 8, 'op': 'literal'}
    instructions[4513] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4514] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4515] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4516] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[4517] = {5'd14, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'unsigned_shift_right'}
    instructions[4518] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4519] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4520] = {5'd1, 4'd8, 4'd4, -32'd2};//{'a': 4, 'literal': -2, 'z': 8, 'op': 'addl'}
    instructions[4521] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[4522] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4523] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4524] = {5'd0, 4'd8, 4'd0, 32'd4};//{'literal': 4, 'z': 8, 'op': 'literal'}
    instructions[4525] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4526] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4527] = {5'd1, 4'd8, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 8, 'op': 'addl'}
    instructions[4528] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4529] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4530] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4531] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[4532] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[4533] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4534] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[4535] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[4536] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4537] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4538] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[4539] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[4540] = {5'd0, 4'd8, 4'd0, 32'd65535};//{'literal': 65535, 'z': 8, 'op': 'literal'}
    instructions[4541] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4542] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4543] = {5'd0, 4'd8, 4'd0, 32'd46};//{'literal': 46, 'z': 8, 'op': 'literal'}
    instructions[4544] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4545] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4546] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4547] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[4548] = {5'd15, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'and'}
    instructions[4549] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4550] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4551] = {5'd1, 4'd8, 4'd4, -32'd2};//{'a': 4, 'literal': -2, 'z': 8, 'op': 'addl'}
    instructions[4552] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[4553] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4554] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4555] = {5'd0, 4'd8, 4'd0, 32'd5};//{'literal': 5, 'z': 8, 'op': 'literal'}
    instructions[4556] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4557] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4558] = {5'd1, 4'd8, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 8, 'op': 'addl'}
    instructions[4559] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4560] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4561] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4562] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[4563] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[4564] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4565] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[4566] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[4567] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4568] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4569] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[4570] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[4571] = {5'd0, 4'd8, 4'd0, 32'd20480};//{'literal': 20480, 'z': 8, 'op': 'literal'}
    instructions[4572] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4573] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4574] = {5'd1, 4'd8, 4'd4, -32'd2};//{'a': 4, 'literal': -2, 'z': 8, 'op': 'addl'}
    instructions[4575] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[4576] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4577] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4578] = {5'd0, 4'd8, 4'd0, 32'd6};//{'literal': 6, 'z': 8, 'op': 'literal'}
    instructions[4579] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4580] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4581] = {5'd1, 4'd8, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 8, 'op': 'addl'}
    instructions[4582] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4583] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4584] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4585] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[4586] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[4587] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4588] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[4589] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[4590] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4591] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4592] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[4593] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[4594] = {5'd0, 4'd8, 4'd0, 32'd1024};//{'literal': 1024, 'z': 8, 'op': 'literal'}
    instructions[4595] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4596] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4597] = {5'd1, 4'd8, 4'd4, -32'd2};//{'a': 4, 'literal': -2, 'z': 8, 'op': 'addl'}
    instructions[4598] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[4599] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4600] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4601] = {5'd0, 4'd8, 4'd0, 32'd7};//{'literal': 7, 'z': 8, 'op': 'literal'}
    instructions[4602] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4603] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4604] = {5'd1, 4'd8, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 8, 'op': 'addl'}
    instructions[4605] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4606] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4607] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4608] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[4609] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[4610] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4611] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[4612] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[4613] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4614] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4615] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[4616] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[4617] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[4618] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4619] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4620] = {5'd1, 4'd8, 4'd4, -32'd2};//{'a': 4, 'literal': -2, 'z': 8, 'op': 'addl'}
    instructions[4621] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[4622] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4623] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4624] = {5'd0, 4'd8, 4'd0, 32'd8};//{'literal': 8, 'z': 8, 'op': 'literal'}
    instructions[4625] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4626] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4627] = {5'd1, 4'd8, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 8, 'op': 'addl'}
    instructions[4628] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4629] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4630] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4631] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[4632] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[4633] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4634] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[4635] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[4636] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4637] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4638] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[4639] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[4640] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[4641] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4642] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4643] = {5'd1, 4'd8, 4'd4, -32'd2};//{'a': 4, 'literal': -2, 'z': 8, 'op': 'addl'}
    instructions[4644] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[4645] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4646] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4647] = {5'd0, 4'd8, 4'd0, 32'd9};//{'literal': 9, 'z': 8, 'op': 'literal'}
    instructions[4648] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4649] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4650] = {5'd1, 4'd8, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 8, 'op': 'addl'}
    instructions[4651] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4652] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4653] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4654] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[4655] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[4656] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4657] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[4658] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[4659] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4660] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4661] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[4662] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[4663] = {5'd0, 4'd8, 4'd0, 32'd2704};//{'literal': 2704, 'z': 8, 'op': 'literal'}
    instructions[4664] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4665] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4666] = {5'd6, 4'd0, 4'd8, 32'd4714};//{'a': 8, 'label': 4714, 'op': 'jmp_if_false'}
    instructions[4667] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[4668] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4669] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4670] = {5'd1, 4'd8, 4'd4, -32'd2};//{'a': 4, 'literal': -2, 'z': 8, 'op': 'addl'}
    instructions[4671] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[4672] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4673] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4674] = {5'd0, 4'd8, 4'd0, 32'd6};//{'literal': 6, 'z': 8, 'op': 'literal'}
    instructions[4675] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4676] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4677] = {5'd1, 4'd8, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 8, 'op': 'addl'}
    instructions[4678] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4679] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4680] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4681] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[4682] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[4683] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4684] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[4685] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[4686] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4687] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4688] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4689] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[4690] = {5'd17, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'or'}
    instructions[4691] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4692] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4693] = {5'd1, 4'd8, 4'd4, -32'd2};//{'a': 4, 'literal': -2, 'z': 8, 'op': 'addl'}
    instructions[4694] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[4695] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4696] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4697] = {5'd0, 4'd8, 4'd0, 32'd6};//{'literal': 6, 'z': 8, 'op': 'literal'}
    instructions[4698] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4699] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4700] = {5'd1, 4'd8, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 8, 'op': 'addl'}
    instructions[4701] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4702] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4703] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4704] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[4705] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[4706] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4707] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[4708] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[4709] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4710] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4711] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[4712] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[4713] = {5'd8, 4'd0, 4'd0, 32'd4714};//{'label': 4714, 'op': 'goto'}
    instructions[4714] = {5'd0, 4'd8, 4'd0, 32'd1079};//{'literal': 1079, 'z': 8, 'op': 'literal'}
    instructions[4715] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4716] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4717] = {5'd6, 4'd0, 4'd8, 32'd4765};//{'a': 8, 'label': 4765, 'op': 'jmp_if_false'}
    instructions[4718] = {5'd0, 4'd8, 4'd0, 32'd2};//{'literal': 2, 'z': 8, 'op': 'literal'}
    instructions[4719] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4720] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4721] = {5'd1, 4'd8, 4'd4, -32'd2};//{'a': 4, 'literal': -2, 'z': 8, 'op': 'addl'}
    instructions[4722] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[4723] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4724] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4725] = {5'd0, 4'd8, 4'd0, 32'd6};//{'literal': 6, 'z': 8, 'op': 'literal'}
    instructions[4726] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4727] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4728] = {5'd1, 4'd8, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 8, 'op': 'addl'}
    instructions[4729] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4730] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4731] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4732] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[4733] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[4734] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4735] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[4736] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[4737] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4738] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4739] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4740] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[4741] = {5'd17, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'or'}
    instructions[4742] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4743] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4744] = {5'd1, 4'd8, 4'd4, -32'd2};//{'a': 4, 'literal': -2, 'z': 8, 'op': 'addl'}
    instructions[4745] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[4746] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4747] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4748] = {5'd0, 4'd8, 4'd0, 32'd6};//{'literal': 6, 'z': 8, 'op': 'literal'}
    instructions[4749] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4750] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4751] = {5'd1, 4'd8, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 8, 'op': 'addl'}
    instructions[4752] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4753] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4754] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4755] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[4756] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[4757] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4758] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[4759] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[4760] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4761] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4762] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[4763] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[4764] = {5'd8, 4'd0, 4'd0, 32'd4765};//{'label': 4765, 'op': 'goto'}
    instructions[4765] = {5'd0, 4'd8, 4'd0, 32'd41};//{'literal': 41, 'z': 8, 'op': 'literal'}
    instructions[4766] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4767] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4768] = {5'd6, 4'd0, 4'd8, 32'd4816};//{'a': 8, 'label': 4816, 'op': 'jmp_if_false'}
    instructions[4769] = {5'd0, 4'd8, 4'd0, 32'd4};//{'literal': 4, 'z': 8, 'op': 'literal'}
    instructions[4770] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4771] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4772] = {5'd1, 4'd8, 4'd4, -32'd2};//{'a': 4, 'literal': -2, 'z': 8, 'op': 'addl'}
    instructions[4773] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[4774] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4775] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4776] = {5'd0, 4'd8, 4'd0, 32'd6};//{'literal': 6, 'z': 8, 'op': 'literal'}
    instructions[4777] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4778] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4779] = {5'd1, 4'd8, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 8, 'op': 'addl'}
    instructions[4780] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4781] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4782] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4783] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[4784] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[4785] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4786] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[4787] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[4788] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4789] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4790] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4791] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[4792] = {5'd17, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'or'}
    instructions[4793] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4794] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4795] = {5'd1, 4'd8, 4'd4, -32'd2};//{'a': 4, 'literal': -2, 'z': 8, 'op': 'addl'}
    instructions[4796] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[4797] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4798] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4799] = {5'd0, 4'd8, 4'd0, 32'd6};//{'literal': 6, 'z': 8, 'op': 'literal'}
    instructions[4800] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4801] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4802] = {5'd1, 4'd8, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 8, 'op': 'addl'}
    instructions[4803] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4804] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4805] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4806] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[4807] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[4808] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4809] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[4810] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[4811] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4812] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4813] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[4814] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[4815] = {5'd8, 4'd0, 4'd0, 32'd4816};//{'label': 4816, 'op': 'goto'}
    instructions[4816] = {5'd0, 4'd8, 4'd0, 32'd34};//{'literal': 34, 'z': 8, 'op': 'literal'}
    instructions[4817] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4818] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4819] = {5'd6, 4'd0, 4'd8, 32'd4867};//{'a': 8, 'label': 4867, 'op': 'jmp_if_false'}
    instructions[4820] = {5'd0, 4'd8, 4'd0, 32'd8};//{'literal': 8, 'z': 8, 'op': 'literal'}
    instructions[4821] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4822] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4823] = {5'd1, 4'd8, 4'd4, -32'd2};//{'a': 4, 'literal': -2, 'z': 8, 'op': 'addl'}
    instructions[4824] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[4825] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4826] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4827] = {5'd0, 4'd8, 4'd0, 32'd6};//{'literal': 6, 'z': 8, 'op': 'literal'}
    instructions[4828] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4829] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4830] = {5'd1, 4'd8, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 8, 'op': 'addl'}
    instructions[4831] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4832] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4833] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4834] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[4835] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[4836] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4837] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[4838] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[4839] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4840] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4841] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4842] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[4843] = {5'd17, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'or'}
    instructions[4844] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4845] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4846] = {5'd1, 4'd8, 4'd4, -32'd2};//{'a': 4, 'literal': -2, 'z': 8, 'op': 'addl'}
    instructions[4847] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[4848] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4849] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4850] = {5'd0, 4'd8, 4'd0, 32'd6};//{'literal': 6, 'z': 8, 'op': 'literal'}
    instructions[4851] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4852] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4853] = {5'd1, 4'd8, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 8, 'op': 'addl'}
    instructions[4854] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4855] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4856] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4857] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[4858] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[4859] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4860] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[4861] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[4862] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4863] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4864] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[4865] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[4866] = {5'd8, 4'd0, 4'd0, 32'd4867};//{'label': 4867, 'op': 'goto'}
    instructions[4867] = {5'd0, 4'd8, 4'd0, 32'd2699};//{'literal': 2699, 'z': 8, 'op': 'literal'}
    instructions[4868] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4869] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4870] = {5'd6, 4'd0, 4'd8, 32'd4918};//{'a': 8, 'label': 4918, 'op': 'jmp_if_false'}
    instructions[4871] = {5'd0, 4'd8, 4'd0, 32'd16};//{'literal': 16, 'z': 8, 'op': 'literal'}
    instructions[4872] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4873] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4874] = {5'd1, 4'd8, 4'd4, -32'd2};//{'a': 4, 'literal': -2, 'z': 8, 'op': 'addl'}
    instructions[4875] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[4876] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4877] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4878] = {5'd0, 4'd8, 4'd0, 32'd6};//{'literal': 6, 'z': 8, 'op': 'literal'}
    instructions[4879] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4880] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4881] = {5'd1, 4'd8, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 8, 'op': 'addl'}
    instructions[4882] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4883] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4884] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4885] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[4886] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[4887] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4888] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[4889] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[4890] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4891] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4892] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4893] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[4894] = {5'd17, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'or'}
    instructions[4895] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4896] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4897] = {5'd1, 4'd8, 4'd4, -32'd2};//{'a': 4, 'literal': -2, 'z': 8, 'op': 'addl'}
    instructions[4898] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[4899] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4900] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4901] = {5'd0, 4'd8, 4'd0, 32'd6};//{'literal': 6, 'z': 8, 'op': 'literal'}
    instructions[4902] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4903] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4904] = {5'd1, 4'd8, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 8, 'op': 'addl'}
    instructions[4905] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4906] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4907] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4908] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[4909] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[4910] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4911] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[4912] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[4913] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4914] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4915] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[4916] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[4917] = {5'd8, 4'd0, 4'd0, 32'd4918};//{'label': 4918, 'op': 'goto'}
    instructions[4918] = {5'd0, 4'd8, 4'd0, 32'd1080};//{'literal': 1080, 'z': 8, 'op': 'literal'}
    instructions[4919] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4920] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4921] = {5'd6, 4'd0, 4'd8, 32'd4969};//{'a': 8, 'label': 4969, 'op': 'jmp_if_false'}
    instructions[4922] = {5'd0, 4'd8, 4'd0, 32'd32};//{'literal': 32, 'z': 8, 'op': 'literal'}
    instructions[4923] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4924] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4925] = {5'd1, 4'd8, 4'd4, -32'd2};//{'a': 4, 'literal': -2, 'z': 8, 'op': 'addl'}
    instructions[4926] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[4927] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4928] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4929] = {5'd0, 4'd8, 4'd0, 32'd6};//{'literal': 6, 'z': 8, 'op': 'literal'}
    instructions[4930] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4931] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4932] = {5'd1, 4'd8, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 8, 'op': 'addl'}
    instructions[4933] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4934] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4935] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4936] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[4937] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[4938] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4939] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[4940] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[4941] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4942] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4943] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4944] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[4945] = {5'd17, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'or'}
    instructions[4946] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4947] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4948] = {5'd1, 4'd8, 4'd4, -32'd2};//{'a': 4, 'literal': -2, 'z': 8, 'op': 'addl'}
    instructions[4949] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[4950] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4951] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4952] = {5'd0, 4'd8, 4'd0, 32'd6};//{'literal': 6, 'z': 8, 'op': 'literal'}
    instructions[4953] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4954] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4955] = {5'd1, 4'd8, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 8, 'op': 'addl'}
    instructions[4956] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4957] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[4958] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4959] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[4960] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[4961] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4962] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[4963] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[4964] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[4965] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4966] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[4967] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[4968] = {5'd8, 4'd0, 4'd0, 32'd4969};//{'label': 4969, 'op': 'goto'}
    instructions[4969] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[4970] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4971] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[4972] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4973] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[4974] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[4975] = {5'd3, 4'd6, 4'd0, 32'd3258};//{'z': 6, 'label': 3258, 'op': 'call'}
    instructions[4976] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[4977] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4978] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[4979] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4980] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[4981] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[4982] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[4983] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4984] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[4985] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4986] = {5'd0, 4'd8, 4'd0, 32'd49320};//{'literal': 49320, 'z': 8, 'op': 'literal'}
    instructions[4987] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[4988] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[4989] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[4990] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[4991] = {5'd3, 4'd6, 4'd0, 32'd3268};//{'z': 6, 'label': 3268, 'op': 'call'}
    instructions[4992] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4993] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4994] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[4995] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[4996] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[4997] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[4998] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[4999] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5000] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[5001] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5002] = {5'd0, 4'd8, 4'd0, 32'd257};//{'literal': 257, 'z': 8, 'op': 'literal'}
    instructions[5003] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5004] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5005] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[5006] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[5007] = {5'd3, 4'd6, 4'd0, 32'd3268};//{'z': 6, 'label': 3268, 'op': 'call'}
    instructions[5008] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5009] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5010] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[5011] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5012] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[5013] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[5014] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[5015] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5016] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[5017] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5018] = {5'd0, 4'd8, 4'd0, 32'd45};//{'literal': 45, 'z': 8, 'op': 'literal'}
    instructions[5019] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5020] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5021] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5022] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5023] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[5024] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[5025] = {5'd3, 4'd6, 4'd0, 32'd3268};//{'z': 6, 'label': 3268, 'op': 'call'}
    instructions[5026] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5027] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5028] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[5029] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5030] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[5031] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[5032] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[5033] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5034] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[5035] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5036] = {5'd0, 4'd8, 4'd0, 32'd1126};//{'literal': 1126, 'z': 8, 'op': 'literal'}
    instructions[5037] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5038] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5039] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5040] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5041] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[5042] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[5043] = {5'd3, 4'd6, 4'd0, 32'd3268};//{'z': 6, 'label': 3268, 'op': 'call'}
    instructions[5044] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5045] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5046] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[5047] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5048] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[5049] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[5050] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[5051] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5052] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[5053] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5054] = {5'd0, 4'd8, 4'd0, 32'd6};//{'literal': 6, 'z': 8, 'op': 'literal'}
    instructions[5055] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5056] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5057] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[5058] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[5059] = {5'd3, 4'd6, 4'd0, 32'd3268};//{'z': 6, 'label': 3268, 'op': 'call'}
    instructions[5060] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5061] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5062] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[5063] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5064] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[5065] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[5066] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[5067] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5068] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[5069] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5070] = {5'd0, 4'd8, 4'd0, 32'd20};//{'literal': 20, 'z': 8, 'op': 'literal'}
    instructions[5071] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5072] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5073] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[5074] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5075] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5076] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5077] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[5078] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[5079] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5080] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5081] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[5082] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[5083] = {5'd3, 4'd6, 4'd0, 32'd3268};//{'z': 6, 'label': 3268, 'op': 'call'}
    instructions[5084] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5085] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5086] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[5087] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5088] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[5089] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[5090] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[5091] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5092] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5093] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[5094] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5095] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5096] = {5'd0, 4'd8, 4'd0, 32'd20};//{'literal': 20, 'z': 8, 'op': 'literal'}
    instructions[5097] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5098] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5099] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[5100] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5101] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5102] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5103] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[5104] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[5105] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5106] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[5107] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[5108] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5109] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[5110] = {5'd14, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'unsigned_shift_right'}
    instructions[5111] = {5'd1, 4'd2, 4'd4, 32'd1};//{'a': 4, 'literal': 1, 'z': 2, 'op': 'addl'}
    instructions[5112] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5113] = {5'd1, 4'd8, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 8, 'op': 'addl'}
    instructions[5114] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5115] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5116] = {5'd1, 4'd2, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 2, 'op': 'addl'}
    instructions[5117] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5118] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[5119] = {5'd1, 4'd2, 4'd4, 32'd3};//{'a': 4, 'literal': 3, 'z': 2, 'op': 'addl'}
    instructions[5120] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5121] = {5'd1, 4'd8, 4'd4, 32'd3};//{'a': 4, 'literal': 3, 'z': 8, 'op': 'addl'}
    instructions[5122] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5123] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5124] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5125] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5126] = {5'd1, 4'd8, 4'd4, 32'd1};//{'a': 4, 'literal': 1, 'z': 8, 'op': 'addl'}
    instructions[5127] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5128] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5129] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5130] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[5131] = {5'd20, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'unsigned_greater'}
    instructions[5132] = {5'd6, 4'd0, 4'd8, 32'd5197};//{'a': 8, 'label': 5197, 'op': 'jmp_if_false'}
    instructions[5133] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[5134] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5135] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[5136] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5137] = {5'd1, 4'd8, 4'd4, -32'd2};//{'a': 4, 'literal': -2, 'z': 8, 'op': 'addl'}
    instructions[5138] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[5139] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5140] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5141] = {5'd1, 4'd8, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 8, 'op': 'addl'}
    instructions[5142] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5143] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5144] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5145] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[5146] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[5147] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5148] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5149] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5150] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5151] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[5152] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[5153] = {5'd3, 4'd6, 4'd0, 32'd3268};//{'z': 6, 'label': 3268, 'op': 'call'}
    instructions[5154] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5155] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5156] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[5157] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5158] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[5159] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[5160] = {5'd1, 4'd8, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 8, 'op': 'addl'}
    instructions[5161] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5162] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5163] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5164] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5165] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[5166] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5167] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5168] = {5'd1, 4'd8, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 8, 'op': 'addl'}
    instructions[5169] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5170] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5171] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5172] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[5173] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[5174] = {5'd1, 4'd2, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 2, 'op': 'addl'}
    instructions[5175] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5176] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5177] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[5178] = {5'd1, 4'd8, 4'd4, 32'd3};//{'a': 4, 'literal': 3, 'z': 8, 'op': 'addl'}
    instructions[5179] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5180] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5181] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5182] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5183] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[5184] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5185] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5186] = {5'd1, 4'd8, 4'd4, 32'd3};//{'a': 4, 'literal': 3, 'z': 8, 'op': 'addl'}
    instructions[5187] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5188] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5189] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5190] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[5191] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[5192] = {5'd1, 4'd2, 4'd4, 32'd3};//{'a': 4, 'literal': 3, 'z': 2, 'op': 'addl'}
    instructions[5193] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5194] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5195] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[5196] = {5'd8, 4'd0, 4'd0, 32'd5121};//{'label': 5121, 'op': 'goto'}
    instructions[5197] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[5198] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5199] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[5200] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5201] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[5202] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[5203] = {5'd3, 4'd6, 4'd0, 32'd3357};//{'z': 6, 'label': 3357, 'op': 'call'}
    instructions[5204] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[5205] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5206] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[5207] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5208] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[5209] = {5'd0, 4'd2, 4'd0, 32'd43};//{'literal': 43, 'z': 2, 'op': 'literal'}
    instructions[5210] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5211] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5212] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5213] = {5'd1, 4'd8, 4'd4, -32'd2};//{'a': 4, 'literal': -2, 'z': 8, 'op': 'addl'}
    instructions[5214] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[5215] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5216] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5217] = {5'd0, 4'd8, 4'd0, 32'd8};//{'literal': 8, 'z': 8, 'op': 'literal'}
    instructions[5218] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5219] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5220] = {5'd1, 4'd8, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 8, 'op': 'addl'}
    instructions[5221] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5222] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5223] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5224] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[5225] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[5226] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5227] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[5228] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[5229] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5230] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5231] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[5232] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5233] = {5'd2, 4'd0, 4'd3, 32'd6};//{'a': 3, 'comment': 'push', 'b': 6, 'op': 'store'}
    instructions[5234] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5235] = {5'd2, 4'd0, 4'd3, 32'd7};//{'a': 3, 'comment': 'push', 'b': 7, 'op': 'store'}
    instructions[5236] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5237] = {5'd1, 4'd8, 4'd4, -32'd2};//{'a': 4, 'literal': -2, 'z': 8, 'op': 'addl'}
    instructions[5238] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[5239] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5240] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5241] = {5'd0, 4'd8, 4'd0, 32'd40};//{'literal': 40, 'z': 8, 'op': 'literal'}
    instructions[5242] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5243] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5244] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[5245] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5246] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5247] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5248] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[5249] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[5250] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5251] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5252] = {5'd0, 4'd8, 4'd0, 32'd6};//{'literal': 6, 'z': 8, 'op': 'literal'}
    instructions[5253] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5254] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5255] = {5'd0, 4'd8, 4'd0, 32'd45};//{'literal': 45, 'z': 8, 'op': 'literal'}
    instructions[5256] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5257] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5258] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5259] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5260] = {5'd0, 4'd8, 4'd0, 32'd1126};//{'literal': 1126, 'z': 8, 'op': 'literal'}
    instructions[5261] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5262] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5263] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5264] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5265] = {5'd1, 4'd7, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 7, 'op': 'addl'}
    instructions[5266] = {5'd1, 4'd4, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[5267] = {5'd3, 4'd6, 4'd0, 32'd3370};//{'z': 6, 'label': 3370, 'op': 'call'}
    instructions[5268] = {5'd1, 4'd3, 4'd3, -32'd5};//{'a': 3, 'literal': -5, 'z': 3, 'op': 'addl'}
    instructions[5269] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5270] = {5'd5, 4'd7, 4'd3, 32'd0};//{'a': 3, 'z': 7, 'op': 'load'}
    instructions[5271] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5272] = {5'd5, 4'd6, 4'd3, 32'd0};//{'a': 3, 'z': 6, 'op': 'load'}
    instructions[5273] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[5274] = {5'd1, 4'd3, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[5275] = {5'd1, 4'd4, 4'd7, 32'd0};//{'a': 7, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[5276] = {5'd12, 4'd0, 4'd6, 32'd0};//{'a': 6, 'op': 'return'}
    instructions[5277] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[5278] = {5'd0, 4'd8, 4'd0, 32'd49};//{'literal': 49, 'z': 8, 'op': 'literal'}
    instructions[5279] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5280] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5281] = {5'd26, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'output_ready'}
    instructions[5282] = {5'd6, 4'd0, 4'd8, 32'd5286};//{'a': 8, 'label': 5286, 'op': 'jmp_if_false'}
    instructions[5283] = {5'd0, 4'd8, 4'd0, 32'd2721};//{'literal': 2721, 'z': 8, 'op': 'literal'}
    instructions[5284] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5285] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5286] = {5'd27, 4'd0, 4'd8, 32'd5301};//{'a': 8, 'label': 5301, 'op': 'jmp_if_true'}
    instructions[5287] = {5'd0, 4'd8, 4'd0, 32'd2154};//{'literal': 2154, 'z': 8, 'op': 'literal'}
    instructions[5288] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5289] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5290] = {5'd21, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'ready'}
    instructions[5291] = {5'd6, 4'd0, 4'd8, 32'd5301};//{'a': 8, 'label': 5301, 'op': 'jmp_if_false'}
    instructions[5292] = {5'd0, 4'd8, 4'd0, 32'd2727};//{'literal': 2727, 'z': 8, 'op': 'literal'}
    instructions[5293] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5294] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5295] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5296] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5297] = {5'd0, 4'd8, 4'd0, 32'd1024};//{'literal': 1024, 'z': 8, 'op': 'literal'}
    instructions[5298] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5299] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[5300] = {5'd19, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'unsigned_greater_equal'}
    instructions[5301] = {5'd6, 4'd0, 4'd8, 32'd5462};//{'a': 8, 'label': 5462, 'op': 'jmp_if_false'}
    instructions[5302] = {5'd0, 4'd8, 4'd0, 32'd49};//{'literal': 49, 'z': 8, 'op': 'literal'}
    instructions[5303] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5304] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5305] = {5'd26, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'output_ready'}
    instructions[5306] = {5'd6, 4'd0, 4'd8, 32'd5310};//{'a': 8, 'label': 5310, 'op': 'jmp_if_false'}
    instructions[5307] = {5'd0, 4'd8, 4'd0, 32'd2721};//{'literal': 2721, 'z': 8, 'op': 'literal'}
    instructions[5308] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5309] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5310] = {5'd6, 4'd0, 4'd8, 32'd5379};//{'a': 8, 'label': 5379, 'op': 'jmp_if_false'}
    instructions[5311] = {5'd0, 4'd8, 4'd0, 32'd49};//{'literal': 49, 'z': 8, 'op': 'literal'}
    instructions[5312] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5313] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5314] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5315] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5316] = {5'd0, 4'd8, 4'd0, 32'd54};//{'literal': 54, 'z': 8, 'op': 'literal'}
    instructions[5317] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5318] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5319] = {5'd0, 4'd8, 4'd0, 32'd1123};//{'literal': 1123, 'z': 8, 'op': 'literal'}
    instructions[5320] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5321] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5322] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5323] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5324] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[5325] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5326] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5327] = {5'd0, 4'd8, 4'd0, 32'd1123};//{'literal': 1123, 'z': 8, 'op': 'literal'}
    instructions[5328] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5329] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5330] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5331] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[5332] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[5333] = {5'd0, 4'd2, 4'd0, 32'd1123};//{'literal': 1123, 'z': 2, 'op': 'literal'}
    instructions[5334] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5335] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5336] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[5337] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5338] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[5339] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[5340] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5341] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5342] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5343] = {5'd5, 4'd0, 4'd3, 32'd0};//{'a': 3, 'z': 0, 'op': 'load'}
    instructions[5344] = {5'd13, 4'd0, 4'd0, 32'd8};//{'a': 0, 'b': 8, 'op': 'write'}
    instructions[5345] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[5346] = {5'd0, 4'd8, 4'd0, 32'd2721};//{'literal': 2721, 'z': 8, 'op': 'literal'}
    instructions[5347] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5348] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5349] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5350] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5351] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[5352] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5353] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5354] = {5'd0, 4'd8, 4'd0, 32'd2721};//{'literal': 2721, 'z': 8, 'op': 'literal'}
    instructions[5355] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5356] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5357] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5358] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[5359] = {5'd10, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'subtract'}
    instructions[5360] = {5'd0, 4'd2, 4'd0, 32'd2721};//{'literal': 2721, 'z': 2, 'op': 'literal'}
    instructions[5361] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5362] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5363] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[5364] = {5'd0, 4'd8, 4'd0, 32'd1024};//{'literal': 1024, 'z': 8, 'op': 'literal'}
    instructions[5365] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5366] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5367] = {5'd0, 4'd8, 4'd0, 32'd1123};//{'literal': 1123, 'z': 8, 'op': 'literal'}
    instructions[5368] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5369] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5370] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5371] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[5372] = {5'd7, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'equal'}
    instructions[5373] = {5'd6, 4'd0, 4'd8, 32'd5378};//{'a': 8, 'label': 5378, 'op': 'jmp_if_false'}
    instructions[5374] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[5375] = {5'd0, 4'd2, 4'd0, 32'd1123};//{'literal': 1123, 'z': 2, 'op': 'literal'}
    instructions[5376] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5377] = {5'd8, 4'd0, 4'd0, 32'd5378};//{'label': 5378, 'op': 'goto'}
    instructions[5378] = {5'd8, 4'd0, 4'd0, 32'd5379};//{'label': 5379, 'op': 'goto'}
    instructions[5379] = {5'd0, 4'd8, 4'd0, 32'd2154};//{'literal': 2154, 'z': 8, 'op': 'literal'}
    instructions[5380] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5381] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5382] = {5'd21, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'ready'}
    instructions[5383] = {5'd6, 4'd0, 4'd8, 32'd5393};//{'a': 8, 'label': 5393, 'op': 'jmp_if_false'}
    instructions[5384] = {5'd0, 4'd8, 4'd0, 32'd2727};//{'literal': 2727, 'z': 8, 'op': 'literal'}
    instructions[5385] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5386] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5387] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5388] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5389] = {5'd0, 4'd8, 4'd0, 32'd1024};//{'literal': 1024, 'z': 8, 'op': 'literal'}
    instructions[5390] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5391] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[5392] = {5'd19, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'unsigned_greater_equal'}
    instructions[5393] = {5'd6, 4'd0, 4'd8, 32'd5461};//{'a': 8, 'label': 5461, 'op': 'jmp_if_false'}
    instructions[5394] = {5'd0, 4'd8, 4'd0, 32'd2154};//{'literal': 2154, 'z': 8, 'op': 'literal'}
    instructions[5395] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5396] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5397] = {5'd22, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'read'}
    instructions[5398] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5399] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5400] = {5'd0, 4'd8, 4'd0, 32'd1130};//{'literal': 1130, 'z': 8, 'op': 'literal'}
    instructions[5401] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5402] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5403] = {5'd0, 4'd8, 4'd0, 32'd53};//{'literal': 53, 'z': 8, 'op': 'literal'}
    instructions[5404] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5405] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5406] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5407] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5408] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[5409] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5410] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5411] = {5'd0, 4'd8, 4'd0, 32'd53};//{'literal': 53, 'z': 8, 'op': 'literal'}
    instructions[5412] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5413] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5414] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5415] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[5416] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[5417] = {5'd0, 4'd2, 4'd0, 32'd53};//{'literal': 53, 'z': 2, 'op': 'literal'}
    instructions[5418] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5419] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5420] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[5421] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5422] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[5423] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[5424] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5425] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5426] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[5427] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5428] = {5'd0, 4'd8, 4'd0, 32'd2727};//{'literal': 2727, 'z': 8, 'op': 'literal'}
    instructions[5429] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5430] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5431] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5432] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5433] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[5434] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5435] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5436] = {5'd0, 4'd8, 4'd0, 32'd2727};//{'literal': 2727, 'z': 8, 'op': 'literal'}
    instructions[5437] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5438] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5439] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5440] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[5441] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[5442] = {5'd0, 4'd2, 4'd0, 32'd2727};//{'literal': 2727, 'z': 2, 'op': 'literal'}
    instructions[5443] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5444] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5445] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[5446] = {5'd0, 4'd8, 4'd0, 32'd1024};//{'literal': 1024, 'z': 8, 'op': 'literal'}
    instructions[5447] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5448] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5449] = {5'd0, 4'd8, 4'd0, 32'd53};//{'literal': 53, 'z': 8, 'op': 'literal'}
    instructions[5450] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5451] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5452] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5453] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[5454] = {5'd7, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'equal'}
    instructions[5455] = {5'd6, 4'd0, 4'd8, 32'd5460};//{'a': 8, 'label': 5460, 'op': 'jmp_if_false'}
    instructions[5456] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[5457] = {5'd0, 4'd2, 4'd0, 32'd53};//{'literal': 53, 'z': 2, 'op': 'literal'}
    instructions[5458] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5459] = {5'd8, 4'd0, 4'd0, 32'd5460};//{'label': 5460, 'op': 'goto'}
    instructions[5460] = {5'd8, 4'd0, 4'd0, 32'd5461};//{'label': 5461, 'op': 'goto'}
    instructions[5461] = {5'd8, 4'd0, 4'd0, 32'd5463};//{'label': 5463, 'op': 'goto'}
    instructions[5462] = {5'd8, 4'd0, 4'd0, 32'd5464};//{'label': 5464, 'op': 'goto'}
    instructions[5463] = {5'd8, 4'd0, 4'd0, 32'd5278};//{'label': 5278, 'op': 'goto'}
    instructions[5464] = {5'd1, 4'd3, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[5465] = {5'd1, 4'd4, 4'd7, 32'd0};//{'a': 7, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[5466] = {5'd12, 4'd0, 4'd6, 32'd0};//{'a': 6, 'op': 'return'}
    instructions[5467] = {5'd1, 4'd3, 4'd3, 32'd6};//{'a': 3, 'literal': 6, 'z': 3, 'op': 'addl'}
    instructions[5468] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[5469] = {5'd1, 4'd2, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5470] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5471] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[5472] = {5'd1, 4'd2, 4'd4, 32'd1};//{'a': 4, 'literal': 1, 'z': 2, 'op': 'addl'}
    instructions[5473] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5474] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[5475] = {5'd1, 4'd2, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 2, 'op': 'addl'}
    instructions[5476] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5477] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[5478] = {5'd1, 4'd2, 4'd4, 32'd3};//{'a': 4, 'literal': 3, 'z': 2, 'op': 'addl'}
    instructions[5479] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5480] = {5'd0, 4'd8, 4'd0, 32'd1090};//{'literal': 1090, 'z': 8, 'op': 'literal'}
    instructions[5481] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5482] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5483] = {5'd1, 4'd2, 4'd4, 32'd4};//{'a': 4, 'literal': 4, 'z': 2, 'op': 'addl'}
    instructions[5484] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5485] = {5'd0, 4'd8, 4'd0, 32'd2727};//{'literal': 2727, 'z': 8, 'op': 'literal'}
    instructions[5486] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5487] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5488] = {5'd1, 4'd2, 4'd4, 32'd5};//{'a': 4, 'literal': 5, 'z': 2, 'op': 'addl'}
    instructions[5489] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5490] = {5'd1, 4'd8, 4'd4, 32'd5};//{'a': 4, 'literal': 5, 'z': 8, 'op': 'addl'}
    instructions[5491] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5492] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5493] = {5'd6, 4'd0, 4'd8, 32'd5711};//{'a': 8, 'label': 5711, 'op': 'jmp_if_false'}
    instructions[5494] = {5'd1, 4'd8, 4'd4, 32'd1};//{'a': 4, 'literal': 1, 'z': 8, 'op': 'addl'}
    instructions[5495] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5496] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5497] = {5'd6, 4'd0, 4'd8, 32'd5558};//{'a': 8, 'label': 5558, 'op': 'jmp_if_false'}
    instructions[5498] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[5499] = {5'd1, 4'd2, 4'd4, 32'd1};//{'a': 4, 'literal': 1, 'z': 2, 'op': 'addl'}
    instructions[5500] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5501] = {5'd0, 4'd8, 4'd0, 32'd8};//{'literal': 8, 'z': 8, 'op': 'literal'}
    instructions[5502] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5503] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5504] = {5'd0, 4'd8, 4'd0, 32'd1130};//{'literal': 1130, 'z': 8, 'op': 'literal'}
    instructions[5505] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5506] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5507] = {5'd1, 4'd8, 4'd4, 32'd4};//{'a': 4, 'literal': 4, 'z': 8, 'op': 'addl'}
    instructions[5508] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5509] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5510] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5511] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5512] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[5513] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5514] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5515] = {5'd1, 4'd8, 4'd4, 32'd4};//{'a': 4, 'literal': 4, 'z': 8, 'op': 'addl'}
    instructions[5516] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5517] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5518] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5519] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[5520] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[5521] = {5'd1, 4'd2, 4'd4, 32'd4};//{'a': 4, 'literal': 4, 'z': 2, 'op': 'addl'}
    instructions[5522] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5523] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5524] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[5525] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5526] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[5527] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[5528] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5529] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5530] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5531] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[5532] = {5'd16, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'shift_left'}
    instructions[5533] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5534] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5535] = {5'd1, 4'd8, 4'd4, -32'd2};//{'a': 4, 'literal': -2, 'z': 8, 'op': 'addl'}
    instructions[5536] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[5537] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5538] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5539] = {5'd1, 4'd8, 4'd4, 32'd3};//{'a': 4, 'literal': 3, 'z': 8, 'op': 'addl'}
    instructions[5540] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5541] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5542] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5543] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5544] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[5545] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5546] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5547] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5548] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[5549] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[5550] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5551] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[5552] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[5553] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5554] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5555] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[5556] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5557] = {5'd8, 4'd0, 4'd0, 32'd5660};//{'label': 5660, 'op': 'goto'}
    instructions[5558] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[5559] = {5'd1, 4'd2, 4'd4, 32'd1};//{'a': 4, 'literal': 1, 'z': 2, 'op': 'addl'}
    instructions[5560] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5561] = {5'd0, 4'd8, 4'd0, 32'd255};//{'literal': 255, 'z': 8, 'op': 'literal'}
    instructions[5562] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5563] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5564] = {5'd0, 4'd8, 4'd0, 32'd1130};//{'literal': 1130, 'z': 8, 'op': 'literal'}
    instructions[5565] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5566] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5567] = {5'd1, 4'd8, 4'd4, 32'd4};//{'a': 4, 'literal': 4, 'z': 8, 'op': 'addl'}
    instructions[5568] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5569] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5570] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5571] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5572] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[5573] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5574] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5575] = {5'd1, 4'd8, 4'd4, 32'd4};//{'a': 4, 'literal': 4, 'z': 8, 'op': 'addl'}
    instructions[5576] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5577] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5578] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5579] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[5580] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[5581] = {5'd1, 4'd2, 4'd4, 32'd4};//{'a': 4, 'literal': 4, 'z': 2, 'op': 'addl'}
    instructions[5582] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5583] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5584] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[5585] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5586] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[5587] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[5588] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5589] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5590] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5591] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[5592] = {5'd15, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'and'}
    instructions[5593] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5594] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5595] = {5'd1, 4'd8, 4'd4, -32'd2};//{'a': 4, 'literal': -2, 'z': 8, 'op': 'addl'}
    instructions[5596] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[5597] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5598] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5599] = {5'd1, 4'd8, 4'd4, 32'd3};//{'a': 4, 'literal': 3, 'z': 8, 'op': 'addl'}
    instructions[5600] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5601] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5602] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5603] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5604] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[5605] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5606] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5607] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5608] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[5609] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[5610] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5611] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[5612] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[5613] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5614] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5615] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5616] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[5617] = {5'd17, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'or'}
    instructions[5618] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5619] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5620] = {5'd1, 4'd8, 4'd4, -32'd2};//{'a': 4, 'literal': -2, 'z': 8, 'op': 'addl'}
    instructions[5621] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[5622] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5623] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5624] = {5'd1, 4'd8, 4'd4, 32'd3};//{'a': 4, 'literal': 3, 'z': 8, 'op': 'addl'}
    instructions[5625] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5626] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5627] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5628] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5629] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[5630] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5631] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5632] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5633] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[5634] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[5635] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5636] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[5637] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[5638] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5639] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5640] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[5641] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5642] = {5'd1, 4'd8, 4'd4, 32'd3};//{'a': 4, 'literal': 3, 'z': 8, 'op': 'addl'}
    instructions[5643] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5644] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5645] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5646] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5647] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[5648] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5649] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5650] = {5'd1, 4'd8, 4'd4, 32'd3};//{'a': 4, 'literal': 3, 'z': 8, 'op': 'addl'}
    instructions[5651] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5652] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5653] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5654] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[5655] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[5656] = {5'd1, 4'd2, 4'd4, 32'd3};//{'a': 4, 'literal': 3, 'z': 2, 'op': 'addl'}
    instructions[5657] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5658] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5659] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[5660] = {5'd0, 4'd8, 4'd0, 32'd1024};//{'literal': 1024, 'z': 8, 'op': 'literal'}
    instructions[5661] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5662] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5663] = {5'd1, 4'd8, 4'd4, 32'd4};//{'a': 4, 'literal': 4, 'z': 8, 'op': 'addl'}
    instructions[5664] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5665] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5666] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5667] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[5668] = {5'd7, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'equal'}
    instructions[5669] = {5'd6, 4'd0, 4'd8, 32'd5674};//{'a': 8, 'label': 5674, 'op': 'jmp_if_false'}
    instructions[5670] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[5671] = {5'd1, 4'd2, 4'd4, 32'd4};//{'a': 4, 'literal': 4, 'z': 2, 'op': 'addl'}
    instructions[5672] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5673] = {5'd8, 4'd0, 4'd0, 32'd5674};//{'label': 5674, 'op': 'goto'}
    instructions[5674] = {5'd1, 4'd8, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 8, 'op': 'addl'}
    instructions[5675] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5676] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5677] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5678] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5679] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[5680] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5681] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5682] = {5'd1, 4'd8, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 8, 'op': 'addl'}
    instructions[5683] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5684] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5685] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5686] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[5687] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[5688] = {5'd1, 4'd2, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5689] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5690] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5691] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[5692] = {5'd1, 4'd8, 4'd4, 32'd5};//{'a': 4, 'literal': 5, 'z': 8, 'op': 'addl'}
    instructions[5693] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5694] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5695] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5696] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5697] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[5698] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5699] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5700] = {5'd1, 4'd8, 4'd4, 32'd5};//{'a': 4, 'literal': 5, 'z': 8, 'op': 'addl'}
    instructions[5701] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5702] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5703] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5704] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[5705] = {5'd10, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'subtract'}
    instructions[5706] = {5'd1, 4'd2, 4'd4, 32'd5};//{'a': 4, 'literal': 5, 'z': 2, 'op': 'addl'}
    instructions[5707] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5708] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5709] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[5710] = {5'd8, 4'd0, 4'd0, 32'd5712};//{'label': 5712, 'op': 'goto'}
    instructions[5711] = {5'd8, 4'd0, 4'd0, 32'd5713};//{'label': 5713, 'op': 'goto'}
    instructions[5712] = {5'd8, 4'd0, 4'd0, 32'd5490};//{'label': 5490, 'op': 'goto'}
    instructions[5713] = {5'd1, 4'd8, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 8, 'op': 'addl'}
    instructions[5714] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5715] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5716] = {5'd0, 4'd2, 4'd0, 32'd2155};//{'literal': 2155, 'z': 2, 'op': 'literal'}
    instructions[5717] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5718] = {5'd1, 4'd3, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[5719] = {5'd1, 4'd4, 4'd7, 32'd0};//{'a': 7, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[5720] = {5'd12, 4'd0, 4'd6, 32'd0};//{'a': 6, 'op': 'return'}
    instructions[5721] = {5'd1, 4'd3, 4'd3, 32'd4};//{'a': 3, 'literal': 4, 'z': 3, 'op': 'addl'}
    instructions[5722] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[5723] = {5'd1, 4'd2, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5724] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5725] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[5726] = {5'd1, 4'd2, 4'd4, 32'd1};//{'a': 4, 'literal': 1, 'z': 2, 'op': 'addl'}
    instructions[5727] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5728] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[5729] = {5'd1, 4'd2, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 2, 'op': 'addl'}
    instructions[5730] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5731] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[5732] = {5'd1, 4'd2, 4'd4, 32'd3};//{'a': 4, 'literal': 3, 'z': 2, 'op': 'addl'}
    instructions[5733] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5734] = {5'd0, 4'd8, 4'd0, 32'd2721};//{'literal': 2721, 'z': 8, 'op': 'literal'}
    instructions[5735] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5736] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5737] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5738] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5739] = {5'd0, 4'd8, 4'd0, 32'd1024};//{'literal': 1024, 'z': 8, 'op': 'literal'}
    instructions[5740] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5741] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[5742] = {5'd10, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'subtract'}
    instructions[5743] = {5'd1, 4'd2, 4'd4, 32'd1};//{'a': 4, 'literal': 1, 'z': 2, 'op': 'addl'}
    instructions[5744] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5745] = {5'd1, 4'd8, 4'd4, 32'd1};//{'a': 4, 'literal': 1, 'z': 8, 'op': 'addl'}
    instructions[5746] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5747] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5748] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5749] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5750] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[5751] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5752] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5753] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5754] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[5755] = {5'd20, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'unsigned_greater'}
    instructions[5756] = {5'd6, 4'd0, 4'd8, 32'd5764};//{'a': 8, 'label': 5764, 'op': 'jmp_if_false'}
    instructions[5757] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[5758] = {5'd0, 4'd2, 4'd0, 32'd2700};//{'literal': 2700, 'z': 2, 'op': 'literal'}
    instructions[5759] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5760] = {5'd1, 4'd3, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[5761] = {5'd1, 4'd4, 4'd7, 32'd0};//{'a': 7, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[5762] = {5'd12, 4'd0, 4'd6, 32'd0};//{'a': 6, 'op': 'return'}
    instructions[5763] = {5'd8, 4'd0, 4'd0, 32'd5764};//{'label': 5764, 'op': 'goto'}
    instructions[5764] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[5765] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5766] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5767] = {5'd6, 4'd0, 4'd8, 32'd5937};//{'a': 8, 'label': 5937, 'op': 'jmp_if_false'}
    instructions[5768] = {5'd1, 4'd8, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 8, 'op': 'addl'}
    instructions[5769] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5770] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5771] = {5'd6, 4'd0, 4'd8, 32'd5804};//{'a': 8, 'label': 5804, 'op': 'jmp_if_false'}
    instructions[5772] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[5773] = {5'd1, 4'd2, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5774] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5775] = {5'd0, 4'd8, 4'd0, 32'd8};//{'literal': 8, 'z': 8, 'op': 'literal'}
    instructions[5776] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5777] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5778] = {5'd1, 4'd8, 4'd4, -32'd3};//{'a': 4, 'literal': -3, 'z': 8, 'op': 'addl'}
    instructions[5779] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[5780] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5781] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5782] = {5'd1, 4'd8, 4'd4, 32'd3};//{'a': 4, 'literal': 3, 'z': 8, 'op': 'addl'}
    instructions[5783] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5784] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5785] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5786] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5787] = {5'd1, 4'd8, 4'd4, -32'd2};//{'a': 4, 'literal': -2, 'z': 8, 'op': 'addl'}
    instructions[5788] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5789] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5790] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5791] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[5792] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[5793] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5794] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[5795] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[5796] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5797] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5798] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5799] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[5800] = {5'd14, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'unsigned_shift_right'}
    instructions[5801] = {5'd1, 4'd2, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 2, 'op': 'addl'}
    instructions[5802] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5803] = {5'd8, 4'd0, 4'd0, 32'd5853};//{'label': 5853, 'op': 'goto'}
    instructions[5804] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[5805] = {5'd1, 4'd2, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5806] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5807] = {5'd0, 4'd8, 4'd0, 32'd255};//{'literal': 255, 'z': 8, 'op': 'literal'}
    instructions[5808] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5809] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5810] = {5'd1, 4'd8, 4'd4, -32'd3};//{'a': 4, 'literal': -3, 'z': 8, 'op': 'addl'}
    instructions[5811] = {5'd5, 4'd8, 4'd8, 32'd0};//{'a': 8, 'z': 8, 'op': 'load'}
    instructions[5812] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5813] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5814] = {5'd1, 4'd8, 4'd4, 32'd3};//{'a': 4, 'literal': 3, 'z': 8, 'op': 'addl'}
    instructions[5815] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5816] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5817] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5818] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5819] = {5'd1, 4'd8, 4'd4, -32'd2};//{'a': 4, 'literal': -2, 'z': 8, 'op': 'addl'}
    instructions[5820] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5821] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5822] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5823] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[5824] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[5825] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5826] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[5827] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[5828] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5829] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5830] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5831] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[5832] = {5'd15, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'and'}
    instructions[5833] = {5'd1, 4'd2, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 2, 'op': 'addl'}
    instructions[5834] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5835] = {5'd1, 4'd8, 4'd4, 32'd3};//{'a': 4, 'literal': 3, 'z': 8, 'op': 'addl'}
    instructions[5836] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5837] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5838] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5839] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5840] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[5841] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5842] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5843] = {5'd1, 4'd8, 4'd4, 32'd3};//{'a': 4, 'literal': 3, 'z': 8, 'op': 'addl'}
    instructions[5844] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5845] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5846] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5847] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[5848] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[5849] = {5'd1, 4'd2, 4'd4, 32'd3};//{'a': 4, 'literal': 3, 'z': 2, 'op': 'addl'}
    instructions[5850] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5851] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5852] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[5853] = {5'd1, 4'd8, 4'd4, 32'd2};//{'a': 4, 'literal': 2, 'z': 8, 'op': 'addl'}
    instructions[5854] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5855] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5856] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5857] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5858] = {5'd0, 4'd8, 4'd0, 32'd54};//{'literal': 54, 'z': 8, 'op': 'literal'}
    instructions[5859] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5860] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5861] = {5'd0, 4'd8, 4'd0, 32'd16};//{'literal': 16, 'z': 8, 'op': 'literal'}
    instructions[5862] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5863] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5864] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5865] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5866] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[5867] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5868] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5869] = {5'd0, 4'd8, 4'd0, 32'd16};//{'literal': 16, 'z': 8, 'op': 'literal'}
    instructions[5870] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5871] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5872] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5873] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[5874] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[5875] = {5'd0, 4'd2, 4'd0, 32'd16};//{'literal': 16, 'z': 2, 'op': 'literal'}
    instructions[5876] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5877] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5878] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[5879] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5880] = {5'd5, 4'd2, 4'd3, 32'd0};//{'a': 3, 'z': 2, 'op': 'load'}
    instructions[5881] = {5'd9, 4'd8, 4'd8, 32'd2};//{'a': 8, 'z': 8, 'b': 2, 'op': 'add'}
    instructions[5882] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5883] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5884] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[5885] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5886] = {5'd0, 4'd8, 4'd0, 32'd1024};//{'literal': 1024, 'z': 8, 'op': 'literal'}
    instructions[5887] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5888] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5889] = {5'd0, 4'd8, 4'd0, 32'd16};//{'literal': 16, 'z': 8, 'op': 'literal'}
    instructions[5890] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5891] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5892] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5893] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[5894] = {5'd7, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'equal'}
    instructions[5895] = {5'd6, 4'd0, 4'd8, 32'd5900};//{'a': 8, 'label': 5900, 'op': 'jmp_if_false'}
    instructions[5896] = {5'd0, 4'd8, 4'd0, 32'd0};//{'literal': 0, 'z': 8, 'op': 'literal'}
    instructions[5897] = {5'd0, 4'd2, 4'd0, 32'd16};//{'literal': 16, 'z': 2, 'op': 'literal'}
    instructions[5898] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5899] = {5'd8, 4'd0, 4'd0, 32'd5900};//{'label': 5900, 'op': 'goto'}
    instructions[5900] = {5'd0, 4'd8, 4'd0, 32'd2721};//{'literal': 2721, 'z': 8, 'op': 'literal'}
    instructions[5901] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5902] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5903] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5904] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5905] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[5906] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5907] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5908] = {5'd0, 4'd8, 4'd0, 32'd2721};//{'literal': 2721, 'z': 8, 'op': 'literal'}
    instructions[5909] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5910] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5911] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5912] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[5913] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[5914] = {5'd0, 4'd2, 4'd0, 32'd2721};//{'literal': 2721, 'z': 2, 'op': 'literal'}
    instructions[5915] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5916] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5917] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[5918] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[5919] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5920] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5921] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5922] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5923] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[5924] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5925] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5926] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[5927] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5928] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5929] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5930] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[5931] = {5'd10, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'subtract'}
    instructions[5932] = {5'd1, 4'd2, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 2, 'op': 'addl'}
    instructions[5933] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5934] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5935] = {5'd5, 4'd8, 4'd3, 32'd0};//{'a': 3, 'z': 8, 'op': 'load'}
    instructions[5936] = {5'd8, 4'd0, 4'd0, 32'd5938};//{'label': 5938, 'op': 'goto'}
    instructions[5937] = {5'd8, 4'd0, 4'd0, 32'd5939};//{'label': 5939, 'op': 'goto'}
    instructions[5938] = {5'd8, 4'd0, 4'd0, 32'd5764};//{'label': 5764, 'op': 'goto'}
    instructions[5939] = {5'd0, 4'd8, 4'd0, 32'd1};//{'literal': 1, 'z': 8, 'op': 'literal'}
    instructions[5940] = {5'd0, 4'd2, 4'd0, 32'd2700};//{'literal': 2700, 'z': 2, 'op': 'literal'}
    instructions[5941] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5942] = {5'd1, 4'd3, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[5943] = {5'd1, 4'd4, 4'd7, 32'd0};//{'a': 7, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[5944] = {5'd12, 4'd0, 4'd6, 32'd0};//{'a': 6, 'op': 'return'}
    instructions[5945] = {5'd1, 4'd3, 4'd3, 32'd0};//{'a': 3, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[5946] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[5947] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5948] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5949] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5950] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5951] = {5'd0, 4'd8, 4'd0, 32'd1090};//{'literal': 1090, 'z': 8, 'op': 'literal'}
    instructions[5952] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5953] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5954] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5955] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[5956] = {5'd9, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'add'}
    instructions[5957] = {5'd0, 4'd2, 4'd0, 32'd1090};//{'literal': 1090, 'z': 2, 'op': 'literal'}
    instructions[5958] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5959] = {5'd0, 4'd8, 4'd0, 32'd1024};//{'literal': 1024, 'z': 8, 'op': 'literal'}
    instructions[5960] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5961] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5962] = {5'd0, 4'd8, 4'd0, 32'd1090};//{'literal': 1090, 'z': 8, 'op': 'literal'}
    instructions[5963] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5964] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5965] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5966] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[5967] = {5'd20, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'unsigned_greater'}
    instructions[5968] = {5'd6, 4'd0, 4'd8, 32'd5981};//{'a': 8, 'label': 5981, 'op': 'jmp_if_false'}
    instructions[5969] = {5'd0, 4'd8, 4'd0, 32'd1024};//{'literal': 1024, 'z': 8, 'op': 'literal'}
    instructions[5970] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5971] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5972] = {5'd0, 4'd8, 4'd0, 32'd1090};//{'literal': 1090, 'z': 8, 'op': 'literal'}
    instructions[5973] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5974] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5975] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5976] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[5977] = {5'd10, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'subtract'}
    instructions[5978] = {5'd0, 4'd2, 4'd0, 32'd1090};//{'literal': 1090, 'z': 2, 'op': 'literal'}
    instructions[5979] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5980] = {5'd8, 4'd0, 4'd0, 32'd5981};//{'label': 5981, 'op': 'goto'}
    instructions[5981] = {5'd1, 4'd8, 4'd4, -32'd1};//{'a': 4, 'literal': -1, 'z': 8, 'op': 'addl'}
    instructions[5982] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5983] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5984] = {5'd2, 4'd0, 4'd3, 32'd8};//{'a': 3, 'comment': 'push', 'b': 8, 'op': 'store'}
    instructions[5985] = {5'd1, 4'd3, 4'd3, 32'd1};//{'a': 3, 'literal': 1, 'z': 3, 'op': 'addl'}
    instructions[5986] = {5'd0, 4'd8, 4'd0, 32'd2727};//{'literal': 2727, 'z': 8, 'op': 'literal'}
    instructions[5987] = {5'd1, 4'd2, 4'd8, 32'd0};//{'a': 8, 'literal': 0, 'z': 2, 'op': 'addl'}
    instructions[5988] = {5'd5, 4'd8, 4'd2, 32'd0};//{'a': 2, 'z': 8, 'op': 'load'}
    instructions[5989] = {5'd1, 4'd3, 4'd3, -32'd1};//{'a': 3, 'comment': 'pop', 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[5990] = {5'd5, 4'd10, 4'd3, 32'd0};//{'a': 3, 'z': 10, 'op': 'load'}
    instructions[5991] = {5'd10, 4'd8, 4'd8, 32'd10};//{'a': 8, 'z': 8, 'b': 10, 'op': 'subtract'}
    instructions[5992] = {5'd0, 4'd2, 4'd0, 32'd2727};//{'literal': 2727, 'z': 2, 'op': 'literal'}
    instructions[5993] = {5'd2, 4'd0, 4'd2, 32'd8};//{'a': 2, 'b': 8, 'op': 'store'}
    instructions[5994] = {5'd1, 4'd3, 4'd4, 32'd0};//{'a': 4, 'literal': 0, 'z': 3, 'op': 'addl'}
    instructions[5995] = {5'd1, 4'd4, 4'd7, 32'd0};//{'a': 7, 'literal': 0, 'z': 4, 'op': 'addl'}
    instructions[5996] = {5'd12, 4'd0, 4'd6, 32'd0};//{'a': 6, 'op': 'return'}
  end

  
  always @(posedge clk)
  begin
    load_data <= memory[load_address];
    if(store_enable && state == execute) begin
      memory[store_address] <= store_data;
    end
  end


  //////////////////////////////////////////////////////////////////////////////
  // PIPELINE STAGE 1 -- FETCH INSTRUCTION
  //                                                                            
  
  always @(posedge clk)
  begin
    //implement memory for instructions
    if (state == instruction_fetch || state == operand_fetch || state == execute) begin
      instruction <= instructions[program_counter];
      program_counter_1 <= program_counter;
    end
  end

  assign opcode    = instruction[44:40];
  assign address_z = instruction[39:36];
  assign address_a = instruction[35:32];
  assign address_b = instruction[3:0];
  assign literal   = instruction[31:0];

  //////////////////////////////////////////////////////////////////////////////
  // PIPELINE STAGE 2 -- FETCH OPERANDS
  //                                                                            
  
  always @(posedge clk)
  begin
    if (write_enable) begin
      registers[address_z_3] <= result;
    end
    if (state == operand_fetch || state == execute) begin
      opcode_2 <= opcode;
      literal_2 <= literal;
      address_a_2 <= address_a;
      address_b_2 <= address_b;
      address_z_2 <= address_z;
      program_counter_2 <= program_counter_1;
    end
  end
  assign register_a = registers[address_a_2];
  assign register_b = registers[address_b_2];
  assign operand_a = (address_a_2 == address_z_3 && write_enable)?result:register_a;
  assign operand_b = (address_b_2 == address_z_3 && write_enable)?result:register_b;
  assign store_address = operand_a;
  assign load_address = operand_a;
  assign store_data = operand_b;
  assign store_enable = (opcode_2==2);

  //////////////////////////////////////////////////////////////////////////////
  // PIPELINE STAGE 3 -- EXECUTE
  //                                                                            
  
  always @(posedge clk)
  begin

  write_enable <= 0;
  case(state)

    //instruction_fetch
    instruction_fetch: begin
      program_counter <= program_counter + 1;
      state <= operand_fetch;
    end
    //operand_fetch
    operand_fetch: begin
      program_counter <= program_counter + 1;
      state <= execute;
    end
    //execute
    execute: begin
      program_counter <= program_counter + 1;
      address_z_3 <= address_z_2;
      case(opcode_2)

        //literal
        16'd0:
        begin
          result<=literal_2;
          write_enable <= 1;
        end

        //addl
        16'd1:
        begin
          result<=operand_a + literal_2;
          write_enable <= 1;
        end

        //store
        16'd2:
        begin
        end

        //call
        16'd3:
        begin
          result <= program_counter_2 + 1;
          write_enable <= 1;
          program_counter <= literal_2;
          state <= instruction_fetch;
        end

        //stop
        16'd4:
        begin
        state <= stop;
        end

        //load
        16'd5:
        begin
          state <= load;
        end

        //jmp_if_false
        16'd6:
        begin
          if (operand_a == 0) begin
            program_counter <= literal_2;
            state <= instruction_fetch;
          end
        end

        //equal
        16'd7:
        begin
          result <= operand_a == operand_b;
          write_enable <= 1;
        end

        //goto
        16'd8:
        begin
          program_counter <= literal_2;
          state <= instruction_fetch;
        end

        //add
        16'd9:
        begin
          long_result = operand_a + operand_b;
          result <= long_result[31:0];
          carry[0] <= long_result[32];
          write_enable <= 1;
        end

        //subtract
        16'd10:
        begin
          long_result = operand_a + (~operand_b) + 1;
          result <= long_result[31:0];
          carry[0] <= ~long_result[32];
          write_enable <= 1;
        end

        //wait_clocks
        16'd11:
        begin
          timer <= operand_a;
          state <= wait_state;
        end

        //return
        16'd12:
        begin
          program_counter <= operand_a;
          state <= instruction_fetch;
        end

        //write
        16'd13:
        begin
          state <= write;
          write_output <= operand_a;
          write_value <= operand_b;
        end

        //unsigned_shift_right
        16'd14:
        begin
          if(operand_b < 32) begin
            result <= operand_a >> operand_b;
            carry <= operand_a << (32-operand_b);
          end else begin
            result <= 0;
            carry <= operand_a;
          end
          write_enable <= 1;
        end

        //and
        16'd15:
        begin
          result <= operand_a & operand_b;
          write_enable <= 1;
        end

        //shift_left
        16'd16:
        begin
          if(operand_b < 32) begin
            result <= operand_a << operand_b;
            carry <= operand_a >> (32-operand_b);
          end else begin
            result <= 0;
            carry <= operand_a;
          end
          write_enable <= 1;
        end

        //or
        16'd17:
        begin
          result <= operand_a | operand_b;
          write_enable <= 1;
        end

        //not_equal
        16'd18:
        begin
          result <= operand_a != operand_b;
          write_enable <= 1;
        end

        //unsigned_greater_equal
        16'd19:
        begin
          result <= $unsigned(operand_a) >= $unsigned(operand_b);
          write_enable <= 1;
        end

        //unsigned_greater
        16'd20:
        begin
          result <= $unsigned(operand_a) > $unsigned(operand_b);
          write_enable <= 1;
        end

        //ready
        16'd21:
        begin
          result <= 0;
          case(operand_a)

            2:
            begin
              result[0] <= input_eth_rx_stb;
            end
            3:
            begin
              result[0] <= input_socket_stb;
            end
          endcase
          write_enable <= 1;
        end

        //read
        16'd22:
        begin
          state <= read;
          read_input <= operand_a;
        end

        //int_to_long
        16'd23:
        begin
          if(operand_a[31]) begin
            result <= -1;
          end else begin
            result <= 0;
          end
          write_enable <= 1;
        end

        //add_with_carry
        16'd24:
        begin
          long_result = operand_a + operand_b + carry[0];
          result <= long_result[31:0];
          carry[0] <= long_result[32];
          write_enable <= 1;
        end

        //not
        16'd25:
        begin
          result <= ~operand_a;
          write_enable <= 1;
        end

        //output_ready
        16'd26:
        begin
          result <= 0;
          case(operand_a)

            0:
            begin
              result[0] <= output_eth_tx_ack;
            end
            1:
            begin
              result[0] <= output_socket_ack;
            end
            4:
            begin
              result[0] <= output_rs232_tx_ack;
            end
          endcase
          write_enable <= 1;
        end

        //jmp_if_true
        16'd27:
        begin
          if (operand_a != 0) begin
            program_counter <= literal_2;
            state <= instruction_fetch;
          end
        end

      endcase

    end

    read:
    begin
      case(read_input)
      2:
      begin
        s_input_eth_rx_ack <= 1;
        if (s_input_eth_rx_ack && input_eth_rx_stb) begin
          result <= input_eth_rx;
          write_enable <= 1;
          s_input_eth_rx_ack <= 0;
          state <= execute;
        end
      end
      3:
      begin
        s_input_socket_ack <= 1;
        if (s_input_socket_ack && input_socket_stb) begin
          result <= input_socket;
          write_enable <= 1;
          s_input_socket_ack <= 0;
          state <= execute;
        end
      end
      endcase
    end

    write:
    begin
      case(write_output)
      0:
      begin
        s_output_eth_tx_stb <= 1;
        s_output_eth_tx <= write_value;
        if (output_eth_tx_ack && s_output_eth_tx_stb) begin
          s_output_eth_tx_stb <= 0;
          state <= execute;
        end
      end
      1:
      begin
        s_output_socket_stb <= 1;
        s_output_socket <= write_value;
        if (output_socket_ack && s_output_socket_stb) begin
          s_output_socket_stb <= 0;
          state <= execute;
        end
      end
      4:
      begin
        s_output_rs232_tx_stb <= 1;
        s_output_rs232_tx <= write_value;
        if (output_rs232_tx_ack && s_output_rs232_tx_stb) begin
          s_output_rs232_tx_stb <= 0;
          state <= execute;
        end
      end
      endcase
    end

    load:
    begin
        result <= load_data;
        write_enable <= 1;
        state <= execute;
    end

    wait_state:
    begin
      if (timer) begin
        timer <= timer - 1;
      end else begin
        state <= execute;
      end
    end

    stop:
    begin
    end

    endcase

    if (rst == 1'b1) begin
      timer <= 0;
      program_counter <= 0;
      address_z_3 <= 0;
      result <= 0;
      a = 0;
      b = 0;
      z = 0;
      state <= instruction_fetch;
      s_input_eth_rx_ack <= 0;
      s_input_socket_ack <= 0;
      s_output_eth_tx_stb <= 0;
      s_output_socket_stb <= 0;
      s_output_rs232_tx_stb <= 0;
    end
  end
  assign input_eth_rx_ack = s_input_eth_rx_ack;
  assign input_socket_ack = s_input_socket_ack;
  assign output_eth_tx_stb = s_output_eth_tx_stb;
  assign output_eth_tx = s_output_eth_tx;
  assign output_socket_stb = s_output_socket_stb;
  assign output_socket = s_output_socket;
  assign output_rs232_tx_stb = s_output_rs232_tx_stb;
  assign output_rs232_tx = s_output_rs232_tx;

endmodule
