//name : main_0
//input : input_i2c_in:16
//output : output_i2c_out:16
//output : output_rs232_tx:16
//source_file : /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c

///+============================================================================+
///|                                                                            |
///|                     This file was generated by Chips                       |
///|                                                                            |
///|                                  Chips                                     |
///|                                                                            |
///|                      http://github.com/dawsonjon/Chips-2.0                 |
///|                                                                            |
///|                                                             Python powered |
///+============================================================================+
module main_0(input_i2c_in,input_i2c_in_stb,output_i2c_out_ack,output_rs232_tx_ack,clk,rst,output_i2c_out,output_rs232_tx,output_i2c_out_stb,output_rs232_tx_stb,input_i2c_in_ack,exception);
  integer file_count;
  reg [31:0] divider_a;
  reg [31:0] divider_b;
  wire [31:0] divider_z;
  reg divider_a_stb;
  wire divider_a_ack;
  reg divider_b_stb;
  wire divider_b_ack;
  wire divider_z_stb;
  reg divider_z_ack;
  reg [31:0] adder_a;
  reg [31:0] adder_b;
  wire [31:0] adder_z;
  reg adder_a_stb;
  wire adder_a_ack;
  reg adder_b_stb;
  wire adder_b_ack;
  wire adder_z_stb;
  reg adder_z_ack;
  reg [31:0] multiplier_a;
  reg [31:0] multiplier_b;
  wire [31:0] multiplier_z;
  reg multiplier_a_stb;
  wire multiplier_a_ack;
  reg multiplier_b_stb;
  wire multiplier_b_ack;
  wire multiplier_z_stb;
  reg multiplier_z_ack;
  reg [31:0] int_to_float_in;
  wire [31:0] int_to_float_out;
  wire int_to_float_out_stb;
  reg int_to_float_out_ack;
  reg int_to_float_in_stb;
  wire int_to_float_in_ack;
  reg [31:0] float_to_int_in;
  wire [31:0] float_to_int_out;
  wire float_to_int_out_stb;
  reg float_to_int_out_ack;
  reg float_to_int_in_stb;
  wire float_to_int_in_ack;
  parameter  stop = 5'd0,
  instruction_fetch = 5'd1,
  operand_fetch = 5'd2,
  execute = 5'd3,
  load = 5'd4,
  wait_state = 5'd5,
  read = 5'd6,
  write = 5'd7,
  divider_write_a = 5'd8,
  divider_write_b = 5'd9,
  divider_read_z = 5'd10,
  adder_write_a = 5'd11,
  adder_write_b = 5'd12,
  adder_read_z = 5'd13,
  multiplier_write_a = 5'd14,
  multiplier_write_b = 5'd15,
  multiplier_read_z = 5'd16,
  int_to_float_write_a = 5'd17,
  int_to_float_read_z = 5'd18,
  float_to_int_write_a = 5'd19,
  float_to_int_read_z = 5'd20;
  input [31:0] input_i2c_in;
  input input_i2c_in_stb;
  input output_i2c_out_ack;
  input output_rs232_tx_ack;
  input clk;
  input rst;
  output [31:0] output_i2c_out;
  output [31:0] output_rs232_tx;
  output output_i2c_out_stb;
  output output_rs232_tx_stb;
  output input_i2c_in_ack;
  reg [31:0] timer;
  reg [63:0] timer_clock;
  reg [15:0] program_counter;
  reg [15:0] program_counter_1;
  reg [15:0] program_counter_2;
  reg [44:0] instruction;
  reg [4:0] opcode_2;
  reg [3:0] a;
  reg [3:0] b;
  reg [3:0] z;
  reg write_enable;
  reg [3:0] address_a_2;
  reg [3:0] address_b_2;
  reg [3:0] address_z_2;
  reg [3:0] address_z_3;
  reg [31:0] load_data;
  reg [31:0] write_output;
  reg [31:0] write_value;
  reg [31:0] read_input;
  reg [15:0] literal_2;
  reg [31:0] a_hi;
  reg [31:0] b_hi;
  reg [31:0] a_lo;
  reg [31:0] b_lo;
  reg [63:0] long_result;
  reg [31:0] result;
  reg [15:0] address;
  reg [31:0] data_out;
  reg [31:0] data_in;
  reg [31:0] carry;
  reg [31:0] s_output_i2c_out_stb;
  reg [31:0] s_output_rs232_tx_stb;
  reg [31:0] s_output_i2c_out;
  reg [31:0] s_output_rs232_tx;
  reg [31:0] s_input_i2c_in_ack;
  reg [20:0] state;
  output reg exception;
  reg [28:0] instructions [1476:0];
  reg [31:0] memory [4096:0];
  reg [31:0] registers [15:0];
  wire [31:0] operand_a;
  wire [31:0] operand_b;
  wire [31:0] register_a;
  wire [31:0] register_b;
  wire [15:0] literal;
  wire [4:0] opcode;
  wire [3:0] address_a;
  wire [3:0] address_b;
  wire [3:0] address_z;
  wire [15:0] load_address;
  wire [15:0] store_address;
  wire [31:0] store_data;
  wire  store_enable;

  //////////////////////////////////////////////////////////////////////////////
  // Floating Point Arithmetic                                                  
  //                                                                            
  // Generate IEEE 754 single precision divider, adder and multiplier           
  //                                                                            
  divider divider_inst(
    .clk(clk),
    .rst(rst),
    .input_a(divider_a),
    .input_a_stb(divider_a_stb),
    .input_a_ack(divider_a_ack),
    .input_b(divider_b),
    .input_b_stb(divider_b_stb),
    .input_b_ack(divider_b_ack),
    .output_z(divider_z),
    .output_z_stb(divider_z_stb),
    .output_z_ack(divider_z_ack)
  );
  adder adder_inst(
    .clk(clk),
    .rst(rst),
    .input_a(adder_a),
    .input_a_stb(adder_a_stb),
    .input_a_ack(adder_a_ack),
    .input_b(adder_b),
    .input_b_stb(adder_b_stb),
    .input_b_ack(adder_b_ack),
    .output_z(adder_z),
    .output_z_stb(adder_z_stb),
    .output_z_ack(adder_z_ack)
  );
  multiplier multiplier_inst(
    .clk(clk),
    .rst(rst),
    .input_a(multiplier_a),
    .input_a_stb(multiplier_a_stb),
    .input_a_ack(multiplier_a_ack),
    .input_b(multiplier_b),
    .input_b_stb(multiplier_b_stb),
    .input_b_ack(multiplier_b_ack),
    .output_z(multiplier_z),
    .output_z_stb(multiplier_z_stb),
    .output_z_ack(multiplier_z_ack)
  );
  int_to_float int_to_float_inst(
    .clk(clk),
    .rst(rst),
    .input_a(int_to_float_in),
    .input_a_stb(int_to_float_in_stb),
    .input_a_ack(int_to_float_in_ack),
    .output_z(int_to_float_out),
    .output_z_stb(int_to_float_out_stb),
    .output_z_ack(int_to_float_out_ack)
  );
  float_to_int float_to_int_inst(
    .clk(clk),
    .rst(rst),
    .input_a(float_to_int_in),
    .input_a_stb(float_to_int_in_stb),
    .input_a_ack(float_to_int_in_ack),
    .output_z(float_to_int_out),
    .output_z_stb(float_to_int_out_stb),
    .output_z_ack(float_to_int_out_ack)
  );

  //////////////////////////////////////////////////////////////////////////////
  // INSTRUCTION INITIALIZATION                                                 
  //                                                                            
  // Initialise the contents of the instruction memory                          
  //
  // Intruction Set
  // ==============
  // 0 {'literal': True, 'op': 'literal'}
  // 1 {'literal': True, 'op': 'addl'}
  // 2 {'literal': False, 'op': 'store'}
  // 3 {'literal': True, 'op': 'call'}
  // 4 {'literal': False, 'op': 'stop'}
  // 5 {'literal': False, 'op': 'load'}
  // 6 {'literal': True, 'op': 'literal_hi'}
  // 7 {'literal': False, 'op': 'a_lo'}
  // 8 {'literal': False, 'op': 'int_to_float'}
  // 9 {'literal': False, 'op': 'float_multiply'}
  // 10 {'literal': False, 'op': 'wait_clocks'}
  // 11 {'literal': True, 'op': 'goto'}
  // 12 {'literal': False, 'op': 'return'}
  // 13 {'literal': False, 'op': 'add'}
  // 14 {'literal': True, 'op': 'jmp_if_false'}
  // 15 {'literal': False, 'op': 'write'}
  // 16 {'literal': False, 'op': 'timer_low'}
  // 17 {'literal': False, 'op': 'unsigned_greater'}
  // 18 {'literal': False, 'op': 'or'}
  // 19 {'literal': False, 'op': 'shift_left'}
  // 20 {'literal': False, 'op': 'unsigned_shift_right'}
  // 21 {'literal': False, 'op': 'read'}
  // 22 {'literal': False, 'op': 'and'}
  // 23 {'literal': False, 'op': 'float_subtract'}
  // 24 {'literal': False, 'op': 'float_divide'}
  // 25 {'literal': False, 'op': 'float_to_int'}
  // 26 {'literal': False, 'op': 'greater'}
  // 27 {'literal': False, 'op': 'subtract'}
  // 28 {'literal': False, 'op': 'greater_equal'}
  // 29 {'literal': False, 'op': 'equal'}
  // Intructions
  // ===========
  
  initial
  begin
    instructions[0] = {5'd0, 4'd3, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 34 {'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 34, 'op': 'literal'}
    instructions[1] = {5'd0, 4'd4, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 34 {'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 34, 'op': 'literal'}
    instructions[2] = {5'd1, 4'd3, 4'd3, 16'd107};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 34 {'a': 3, 'literal': 107, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 34, 'op': 'addl'}
    instructions[3] = {5'd0, 4'd8, 4'd0, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 10, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[4] = {5'd0, 4'd2, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[5] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'store'}
    instructions[6] = {5'd0, 4'd8, 4'd0, 16'd67};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 67, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[7] = {5'd0, 4'd2, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[8] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'store'}
    instructions[9] = {5'd0, 4'd8, 4'd0, 16'd104};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 104, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[10] = {5'd0, 4'd2, 4'd0, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[11] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'store'}
    instructions[12] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[13] = {5'd0, 4'd2, 4'd0, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 4, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[14] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'store'}
    instructions[15] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[16] = {5'd0, 4'd2, 4'd0, 16'd5};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 5, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[17] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'store'}
    instructions[18] = {5'd0, 4'd8, 4'd0, 16'd115};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 115, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[19] = {5'd0, 4'd2, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 6, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[20] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'store'}
    instructions[21] = {5'd0, 4'd8, 4'd0, 16'd45};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 45, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[22] = {5'd0, 4'd2, 4'd0, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 7, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[23] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'store'}
    instructions[24] = {5'd0, 4'd8, 4'd0, 16'd50};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 50, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[25] = {5'd0, 4'd2, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 8, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[26] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'store'}
    instructions[27] = {5'd0, 4'd8, 4'd0, 16'd46};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 46, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[28] = {5'd0, 4'd2, 4'd0, 16'd9};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 9, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[29] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'store'}
    instructions[30] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[31] = {5'd0, 4'd2, 4'd0, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 10, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[32] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'store'}
    instructions[33] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[34] = {5'd0, 4'd2, 4'd0, 16'd11};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 11, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[35] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'store'}
    instructions[36] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[37] = {5'd0, 4'd2, 4'd0, 16'd12};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 12, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[38] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'store'}
    instructions[39] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[40] = {5'd0, 4'd2, 4'd0, 16'd13};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 13, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[41] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'store'}
    instructions[42] = {5'd0, 4'd8, 4'd0, 16'd109};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 109, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[43] = {5'd0, 4'd2, 4'd0, 16'd14};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 14, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[44] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'store'}
    instructions[45] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[46] = {5'd0, 4'd2, 4'd0, 16'd15};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 15, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[47] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'store'}
    instructions[48] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[49] = {5'd0, 4'd2, 4'd0, 16'd16};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 16, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[50] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'store'}
    instructions[51] = {5'd0, 4'd8, 4'd0, 16'd114};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 114, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[52] = {5'd0, 4'd2, 4'd0, 16'd17};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 17, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[53] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'store'}
    instructions[54] = {5'd0, 4'd8, 4'd0, 16'd97};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 97, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[55] = {5'd0, 4'd2, 4'd0, 16'd18};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 18, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[56] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'store'}
    instructions[57] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[58] = {5'd0, 4'd2, 4'd0, 16'd19};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 19, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[59] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'store'}
    instructions[60] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[61] = {5'd0, 4'd2, 4'd0, 16'd20};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 20, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[62] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'store'}
    instructions[63] = {5'd0, 4'd8, 4'd0, 16'd114};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 114, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[64] = {5'd0, 4'd2, 4'd0, 16'd21};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 21, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[65] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'store'}
    instructions[66] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[67] = {5'd0, 4'd2, 4'd0, 16'd22};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 22, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[68] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'store'}
    instructions[69] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[70] = {5'd0, 4'd2, 4'd0, 16'd23};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 23, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[71] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'store'}
    instructions[72] = {5'd0, 4'd8, 4'd0, 16'd115};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 115, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[73] = {5'd0, 4'd2, 4'd0, 16'd24};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 24, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[74] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'store'}
    instructions[75] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[76] = {5'd0, 4'd2, 4'd0, 16'd25};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 25, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[77] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'store'}
    instructions[78] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[79] = {5'd0, 4'd2, 4'd0, 16'd26};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 26, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[80] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'store'}
    instructions[81] = {5'd0, 4'd8, 4'd0, 16'd115};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 115, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[82] = {5'd0, 4'd2, 4'd0, 16'd27};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 27, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[83] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'store'}
    instructions[84] = {5'd0, 4'd8, 4'd0, 16'd111};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 111, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[85] = {5'd0, 4'd2, 4'd0, 16'd28};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 28, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[86] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'store'}
    instructions[87] = {5'd0, 4'd8, 4'd0, 16'd114};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 114, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[88] = {5'd0, 4'd2, 4'd0, 16'd29};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 29, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[89] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'store'}
    instructions[90] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[91] = {5'd0, 4'd2, 4'd0, 16'd30};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 30, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[92] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'store'}
    instructions[93] = {5'd0, 4'd8, 4'd0, 16'd100};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 100, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[94] = {5'd0, 4'd2, 4'd0, 16'd31};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 31, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[95] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'store'}
    instructions[96] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[97] = {5'd0, 4'd2, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 32, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[98] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'store'}
    instructions[99] = {5'd0, 4'd8, 4'd0, 16'd109};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 109, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[100] = {5'd0, 4'd2, 4'd0, 16'd33};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 33, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[101] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'store'}
    instructions[102] = {5'd0, 4'd8, 4'd0, 16'd111};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 111, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[103] = {5'd0, 4'd2, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 34, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[104] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'store'}
    instructions[105] = {5'd0, 4'd8, 4'd0, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 10, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[106] = {5'd0, 4'd2, 4'd0, 16'd35};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 35, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[107] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'store'}
    instructions[108] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[109] = {5'd0, 4'd2, 4'd0, 16'd36};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 36, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[110] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'store'}
    instructions[111] = {5'd0, 4'd8, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 7 {'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 7, 'op': 'literal'}
    instructions[112] = {5'd0, 4'd2, 4'd0, 16'd38};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 7 {'literal': 38, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 7, 'op': 'literal'}
    instructions[113] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 7 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 7, 'op': 'store'}
    instructions[114] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 5 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 5, 'op': 'literal'}
    instructions[115] = {5'd0, 4'd2, 4'd0, 16'd40};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 5 {'literal': 40, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 5, 'op': 'literal'}
    instructions[116] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 5 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 5, 'op': 'store'}
    instructions[117] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'literal'}
    instructions[118] = {5'd0, 4'd2, 4'd0, 16'd41};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'literal': 41, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'literal'}
    instructions[119] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'store'}
    instructions[120] = {5'd0, 4'd8, 4'd0, 16'd100};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'literal': 100, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'literal'}
    instructions[121] = {5'd0, 4'd2, 4'd0, 16'd42};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'literal': 42, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'literal'}
    instructions[122] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'store'}
    instructions[123] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'literal'}
    instructions[124] = {5'd0, 4'd2, 4'd0, 16'd43};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'literal': 43, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'literal'}
    instructions[125] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'store'}
    instructions[126] = {5'd0, 4'd8, 4'd0, 16'd103};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'literal': 103, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'literal'}
    instructions[127] = {5'd0, 4'd2, 4'd0, 16'd44};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'literal': 44, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'literal'}
    instructions[128] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'store'}
    instructions[129] = {5'd0, 4'd8, 4'd0, 16'd114};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'literal': 114, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'literal'}
    instructions[130] = {5'd0, 4'd2, 4'd0, 16'd45};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'literal': 45, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'literal'}
    instructions[131] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'store'}
    instructions[132] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'literal'}
    instructions[133] = {5'd0, 4'd2, 4'd0, 16'd46};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'literal': 46, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'literal'}
    instructions[134] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'store'}
    instructions[135] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'literal'}
    instructions[136] = {5'd0, 4'd2, 4'd0, 16'd47};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'literal': 47, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'literal'}
    instructions[137] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'store'}
    instructions[138] = {5'd0, 4'd8, 4'd0, 16'd115};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'literal': 115, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'literal'}
    instructions[139] = {5'd0, 4'd2, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'literal': 48, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'literal'}
    instructions[140] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'store'}
    instructions[141] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'literal'}
    instructions[142] = {5'd0, 4'd2, 4'd0, 16'd49};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'literal': 49, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'literal'}
    instructions[143] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'store'}
    instructions[144] = {5'd0, 4'd8, 4'd0, 16'd67};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'literal': 67, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'literal'}
    instructions[145] = {5'd0, 4'd2, 4'd0, 16'd50};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'literal': 50, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'literal'}
    instructions[146] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'store'}
    instructions[147] = {5'd0, 4'd8, 4'd0, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'literal': 10, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'literal'}
    instructions[148] = {5'd0, 4'd2, 4'd0, 16'd51};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'literal': 51, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'literal'}
    instructions[149] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'store'}
    instructions[150] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'literal'}
    instructions[151] = {5'd0, 4'd2, 4'd0, 16'd52};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'literal': 52, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'literal'}
    instructions[152] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'store'}
    instructions[153] = {5'd0, 4'd8, 4'd0, 16'd73};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 73, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[154] = {5'd0, 4'd2, 4'd0, 16'd53};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 53, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[155] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'store'}
    instructions[156] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[157] = {5'd0, 4'd2, 4'd0, 16'd54};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 54, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[158] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'store'}
    instructions[159] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[160] = {5'd0, 4'd2, 4'd0, 16'd55};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 55, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[161] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'store'}
    instructions[162] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[163] = {5'd0, 4'd2, 4'd0, 16'd56};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 56, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[164] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'store'}
    instructions[165] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[166] = {5'd0, 4'd2, 4'd0, 16'd57};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 57, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[167] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'store'}
    instructions[168] = {5'd0, 4'd8, 4'd0, 16'd97};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 97, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[169] = {5'd0, 4'd2, 4'd0, 16'd58};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 58, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[170] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'store'}
    instructions[171] = {5'd0, 4'd8, 4'd0, 16'd108};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 108, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[172] = {5'd0, 4'd2, 4'd0, 16'd59};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 59, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[173] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'store'}
    instructions[174] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[175] = {5'd0, 4'd2, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 60, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[176] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'store'}
    instructions[177] = {5'd0, 4'd8, 4'd0, 16'd115};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 115, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[178] = {5'd0, 4'd2, 4'd0, 16'd61};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 61, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[179] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'store'}
    instructions[180] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[181] = {5'd0, 4'd2, 4'd0, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 62, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[182] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'store'}
    instructions[183] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[184] = {5'd0, 4'd2, 4'd0, 16'd63};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 63, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[185] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'store'}
    instructions[186] = {5'd0, 4'd8, 4'd0, 16'd103};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 103, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[187] = {5'd0, 4'd2, 4'd0, 16'd64};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 64, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[188] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'store'}
    instructions[189] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[190] = {5'd0, 4'd2, 4'd0, 16'd65};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 65, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[191] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'store'}
    instructions[192] = {5'd0, 4'd8, 4'd0, 16'd65};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 65, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[193] = {5'd0, 4'd2, 4'd0, 16'd66};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 66, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[194] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'store'}
    instructions[195] = {5'd0, 4'd8, 4'd0, 16'd68};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 68, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[196] = {5'd0, 4'd2, 4'd0, 16'd67};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 67, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[197] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'store'}
    instructions[198] = {5'd0, 4'd8, 4'd0, 16'd84};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 84, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[199] = {5'd0, 4'd2, 4'd0, 16'd68};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 68, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[200] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'store'}
    instructions[201] = {5'd0, 4'd8, 4'd0, 16'd55};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 55, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[202] = {5'd0, 4'd2, 4'd0, 16'd69};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 69, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[203] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'store'}
    instructions[204] = {5'd0, 4'd8, 4'd0, 16'd52};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 52, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[205] = {5'd0, 4'd2, 4'd0, 16'd70};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 70, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[206] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'store'}
    instructions[207] = {5'd0, 4'd8, 4'd0, 16'd50};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 50, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[208] = {5'd0, 4'd2, 4'd0, 16'd71};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 71, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[209] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'store'}
    instructions[210] = {5'd0, 4'd8, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 48, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[211] = {5'd0, 4'd2, 4'd0, 16'd72};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 72, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[212] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'store'}
    instructions[213] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[214] = {5'd0, 4'd2, 4'd0, 16'd73};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 73, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[215] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'store'}
    instructions[216] = {5'd0, 4'd8, 4'd0, 16'd98};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 98, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[217] = {5'd0, 4'd2, 4'd0, 16'd74};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 74, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[218] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'store'}
    instructions[219] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[220] = {5'd0, 4'd2, 4'd0, 16'd75};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 75, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[221] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'store'}
    instructions[222] = {5'd0, 4'd8, 4'd0, 16'd115};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 115, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[223] = {5'd0, 4'd2, 4'd0, 16'd76};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 76, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[224] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'store'}
    instructions[225] = {5'd0, 4'd8, 4'd0, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 10, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[226] = {5'd0, 4'd2, 4'd0, 16'd77};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 77, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[227] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'store'}
    instructions[228] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[229] = {5'd0, 4'd2, 4'd0, 16'd78};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 78, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[230] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'store'}
    instructions[231] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 5 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 5, 'op': 'literal'}
    instructions[232] = {5'd0, 4'd2, 4'd0, 16'd79};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 5 {'literal': 79, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 5, 'op': 'literal'}
    instructions[233] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 5 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 5, 'op': 'store'}
    instructions[234] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 6 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 6, 'op': 'literal'}
    instructions[235] = {5'd0, 4'd2, 4'd0, 16'd81};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 6 {'literal': 81, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 6, 'op': 'literal'}
    instructions[236] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 6 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 6, 'op': 'store'}
    instructions[237] = {5'd0, 4'd8, 4'd0, 16'd73};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'literal': 73, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'literal'}
    instructions[238] = {5'd0, 4'd2, 4'd0, 16'd83};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'literal': 83, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'literal'}
    instructions[239] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'store'}
    instructions[240] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'literal'}
    instructions[241] = {5'd0, 4'd2, 4'd0, 16'd84};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'literal': 84, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'literal'}
    instructions[242] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'store'}
    instructions[243] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'literal'}
    instructions[244] = {5'd0, 4'd2, 4'd0, 16'd85};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'literal': 85, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'literal'}
    instructions[245] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'store'}
    instructions[246] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'literal'}
    instructions[247] = {5'd0, 4'd2, 4'd0, 16'd86};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'literal': 86, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'literal'}
    instructions[248] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'store'}
    instructions[249] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'literal'}
    instructions[250] = {5'd0, 4'd2, 4'd0, 16'd87};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'literal': 87, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'literal'}
    instructions[251] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'store'}
    instructions[252] = {5'd0, 4'd8, 4'd0, 16'd97};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'literal': 97, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'literal'}
    instructions[253] = {5'd0, 4'd2, 4'd0, 16'd88};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'literal': 88, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'literal'}
    instructions[254] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'store'}
    instructions[255] = {5'd0, 4'd8, 4'd0, 16'd108};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'literal': 108, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'literal'}
    instructions[256] = {5'd0, 4'd2, 4'd0, 16'd89};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'literal': 89, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'literal'}
    instructions[257] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'store'}
    instructions[258] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'literal'}
    instructions[259] = {5'd0, 4'd2, 4'd0, 16'd90};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'literal': 90, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'literal'}
    instructions[260] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'store'}
    instructions[261] = {5'd0, 4'd8, 4'd0, 16'd115};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'literal': 115, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'literal'}
    instructions[262] = {5'd0, 4'd2, 4'd0, 16'd91};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'literal': 91, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'literal'}
    instructions[263] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'store'}
    instructions[264] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'literal'}
    instructions[265] = {5'd0, 4'd2, 4'd0, 16'd92};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'literal': 92, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'literal'}
    instructions[266] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'store'}
    instructions[267] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'literal'}
    instructions[268] = {5'd0, 4'd2, 4'd0, 16'd93};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'literal': 93, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'literal'}
    instructions[269] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'store'}
    instructions[270] = {5'd0, 4'd8, 4'd0, 16'd103};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'literal': 103, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'literal'}
    instructions[271] = {5'd0, 4'd2, 4'd0, 16'd94};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'literal': 94, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'literal'}
    instructions[272] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'store'}
    instructions[273] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'literal'}
    instructions[274] = {5'd0, 4'd2, 4'd0, 16'd95};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'literal': 95, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'literal'}
    instructions[275] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'store'}
    instructions[276] = {5'd0, 4'd8, 4'd0, 16'd73};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'literal': 73, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'literal'}
    instructions[277] = {5'd0, 4'd2, 4'd0, 16'd96};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'literal': 96, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'literal'}
    instructions[278] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'store'}
    instructions[279] = {5'd0, 4'd8, 4'd0, 16'd50};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'literal': 50, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'literal'}
    instructions[280] = {5'd0, 4'd2, 4'd0, 16'd97};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'literal': 97, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'literal'}
    instructions[281] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'store'}
    instructions[282] = {5'd0, 4'd8, 4'd0, 16'd67};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'literal': 67, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'literal'}
    instructions[283] = {5'd0, 4'd2, 4'd0, 16'd98};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'literal': 98, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'literal'}
    instructions[284] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'store'}
    instructions[285] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'literal'}
    instructions[286] = {5'd0, 4'd2, 4'd0, 16'd99};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'literal': 99, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'literal'}
    instructions[287] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'store'}
    instructions[288] = {5'd0, 4'd8, 4'd0, 16'd98};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'literal': 98, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'literal'}
    instructions[289] = {5'd0, 4'd2, 4'd0, 16'd100};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'literal': 100, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'literal'}
    instructions[290] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'store'}
    instructions[291] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'literal'}
    instructions[292] = {5'd0, 4'd2, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'literal': 101, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'literal'}
    instructions[293] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'store'}
    instructions[294] = {5'd0, 4'd8, 4'd0, 16'd115};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'literal': 115, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'literal'}
    instructions[295] = {5'd0, 4'd2, 4'd0, 16'd102};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'literal': 102, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'literal'}
    instructions[296] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'store'}
    instructions[297] = {5'd0, 4'd8, 4'd0, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'literal': 10, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'literal'}
    instructions[298] = {5'd0, 4'd2, 4'd0, 16'd103};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'literal': 103, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'literal'}
    instructions[299] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'store'}
    instructions[300] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'literal'}
    instructions[301] = {5'd0, 4'd2, 4'd0, 16'd104};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'literal': 104, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'literal'}
    instructions[302] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'store'}
    instructions[303] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 34 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 34, 'op': 'addl'}
    instructions[304] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 34 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 34, 'op': 'addl'}
    instructions[305] = {5'd3, 4'd6, 4'd0, 16'd307};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 34 {'z': 6, 'label': 307, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 34, 'op': 'call'}
    instructions[306] = {5'd4, 4'd0, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 34 {'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 34, 'op': 'stop'}
    instructions[307] = {5'd1, 4'd3, 4'd3, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 9 {'a': 3, 'literal': 101, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 9, 'op': 'addl'}
    instructions[308] = {5'd0, 4'd8, 4'd0, 16'd38};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 14 {'literal': 38, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 14, 'op': 'literal'}
    instructions[309] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 14 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 14, 'op': 'addl'}
    instructions[310] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 14 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 14, 'op': 'load'}
    instructions[311] = {5'd0, 4'd2, 4'd0, 16'd79};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 14 {'literal': 79, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 14, 'op': 'literal'}
    instructions[312] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 14 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 14, 'op': 'store'}
    instructions[313] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'store'}
    instructions[314] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'addl'}
    instructions[315] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'store'}
    instructions[316] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'addl'}
    instructions[317] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'literal'}
    instructions[318] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'store'}
    instructions[319] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'addl'}
    instructions[320] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'addl'}
    instructions[321] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'addl'}
    instructions[322] = {5'd3, 4'd6, 4'd0, 16'd479};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'z': 6, 'label': 479, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'call'}
    instructions[323] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'addl'}
    instructions[324] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[325] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'load'}
    instructions[326] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[327] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'load'}
    instructions[328] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 16, 'op': 'addl'}
    instructions[329] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'store'}
    instructions[330] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'addl'}
    instructions[331] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'store'}
    instructions[332] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'addl'}
    instructions[333] = {5'd0, 4'd8, 4'd0, 16'd83};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'literal': 83, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'literal'}
    instructions[334] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'store'}
    instructions[335] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'addl'}
    instructions[336] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'addl'}
    instructions[337] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'addl'}
    instructions[338] = {5'd3, 4'd6, 4'd0, 16'd479};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'z': 6, 'label': 479, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'call'}
    instructions[339] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'addl'}
    instructions[340] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[341] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'load'}
    instructions[342] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[343] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'load'}
    instructions[344] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 19, 'op': 'addl'}
    instructions[345] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20, 'op': 'store'}
    instructions[346] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20, 'op': 'addl'}
    instructions[347] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20, 'op': 'store'}
    instructions[348] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20, 'op': 'addl'}
    instructions[349] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20, 'op': 'addl'}
    instructions[350] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20, 'op': 'store'}
    instructions[351] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20, 'op': 'addl'}
    instructions[352] = {5'd0, 4'd8, 4'd0, 16'd40};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20 {'literal': 40, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20, 'op': 'literal'}
    instructions[353] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20, 'op': 'addl'}
    instructions[354] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20, 'op': 'load'}
    instructions[355] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20, 'op': 'store'}
    instructions[356] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20, 'op': 'addl'}
    instructions[357] = {5'd0, 4'd8, 4'd0, 16'd81};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20 {'literal': 81, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20, 'op': 'literal'}
    instructions[358] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20, 'op': 'addl'}
    instructions[359] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20, 'op': 'load'}
    instructions[360] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20, 'op': 'store'}
    instructions[361] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20, 'op': 'addl'}
    instructions[362] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20, 'op': 'addl'}
    instructions[363] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20, 'op': 'addl'}
    instructions[364] = {5'd3, 4'd6, 4'd0, 16'd570};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20 {'z': 6, 'label': 570, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20, 'op': 'call'}
    instructions[365] = {5'd1, 4'd3, 4'd3, -16'd3};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20 {'a': 3, 'literal': -3, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20, 'op': 'addl'}
    instructions[366] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[367] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20, 'op': 'load'}
    instructions[368] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[369] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20, 'op': 'load'}
    instructions[370] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 20, 'op': 'addl'}
    instructions[371] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'store'}
    instructions[372] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'addl'}
    instructions[373] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'store'}
    instructions[374] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'addl'}
    instructions[375] = {5'd0, 4'd8, 4'd0, 16'd53};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'literal': 53, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'literal'}
    instructions[376] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'store'}
    instructions[377] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'addl'}
    instructions[378] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'addl'}
    instructions[379] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'addl'}
    instructions[380] = {5'd3, 4'd6, 4'd0, 16'd479};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'z': 6, 'label': 479, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'call'}
    instructions[381] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'addl'}
    instructions[382] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[383] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'load'}
    instructions[384] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[385] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'load'}
    instructions[386] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 23, 'op': 'addl'}
    instructions[387] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 24 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 24, 'op': 'store'}
    instructions[388] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 24 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 24, 'op': 'addl'}
    instructions[389] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 24 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 24, 'op': 'store'}
    instructions[390] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 24 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 24, 'op': 'addl'}
    instructions[391] = {5'd1, 4'd8, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 24 {'a': 4, 'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 24, 'op': 'addl'}
    instructions[392] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 24 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 24, 'op': 'store'}
    instructions[393] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 24 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 24, 'op': 'addl'}
    instructions[394] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 24 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 24, 'op': 'addl'}
    instructions[395] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 24 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 24, 'op': 'store'}
    instructions[396] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 24 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 24, 'op': 'addl'}
    instructions[397] = {5'd0, 4'd8, 4'd0, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 24 {'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 24, 'op': 'literal'}
    instructions[398] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 24 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 24, 'op': 'store'}
    instructions[399] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 24 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 24, 'op': 'addl'}
    instructions[400] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 24 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 24, 'op': 'addl'}
    instructions[401] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 24 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 24, 'op': 'addl'}
    instructions[402] = {5'd3, 4'd6, 4'd0, 16'd600};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 24 {'z': 6, 'label': 600, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 24, 'op': 'call'}
    instructions[403] = {5'd1, 4'd3, 4'd3, -16'd3};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 24 {'a': 3, 'literal': -3, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 24, 'op': 'addl'}
    instructions[404] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 24 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 24, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[405] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 24 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 24, 'op': 'load'}
    instructions[406] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 24 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 24, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[407] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 24 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 24, 'op': 'load'}
    instructions[408] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 24 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 24, 'op': 'addl'}
    instructions[409] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 28 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 28, 'op': 'store'}
    instructions[410] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 28 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 28, 'op': 'addl'}
    instructions[411] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 28 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 28, 'op': 'store'}
    instructions[412] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 28 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 28, 'op': 'addl'}
    instructions[413] = {5'd1, 4'd8, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 28 {'a': 4, 'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 28, 'op': 'addl'}
    instructions[414] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 28 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 28, 'op': 'store'}
    instructions[415] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 28 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 28, 'op': 'addl'}
    instructions[416] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 28 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 28, 'op': 'addl'}
    instructions[417] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 28 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 28, 'op': 'addl'}
    instructions[418] = {5'd3, 4'd6, 4'd0, 16'd641};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 28 {'z': 6, 'label': 641, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 28, 'op': 'call'}
    instructions[419] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 28 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 28, 'op': 'addl'}
    instructions[420] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 28 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 28, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[421] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 28 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 28, 'op': 'load'}
    instructions[422] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 28 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 28, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[423] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 28 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 28, 'op': 'load'}
    instructions[424] = {5'd0, 4'd2, 4'd0, 16'd37};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 28 {'literal': 37, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 28, 'op': 'literal'}
    instructions[425] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 28 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 28, 'op': 'load'}
    instructions[426] = {5'd1, 4'd2, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 28 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 28, 'op': 'addl'}
    instructions[427] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 28 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 28, 'op': 'store'}
    instructions[428] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29, 'op': 'store'}
    instructions[429] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29, 'op': 'addl'}
    instructions[430] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29, 'op': 'store'}
    instructions[431] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29, 'op': 'addl'}
    instructions[432] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29, 'op': 'literal'}
    instructions[433] = {5'd6, 4'd8, 4'd8, 16'd15744};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29 {'a': 8, 'literal': 15744, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29, 'op': 'literal_hi'}
    instructions[434] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29, 'op': 'store'}
    instructions[435] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29, 'op': 'addl'}
    instructions[436] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29, 'op': 'addl'}
    instructions[437] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29, 'op': 'addl'}
    instructions[438] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29, 'op': 'load'}
    instructions[439] = {5'd7, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29 {'a': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29, 'op': 'a_lo'}
    instructions[440] = {5'd8, 4'd0, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29 {'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29, 'op': 'int_to_float'}
    instructions[441] = {5'd7, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29 {'a': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29, 'op': 'a_lo'}
    instructions[442] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[443] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29, 'op': 'load'}
    instructions[444] = {5'd9, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29, 'op': 'float_multiply'}
    instructions[445] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29, 'op': 'store'}
    instructions[446] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29, 'op': 'addl'}
    instructions[447] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29, 'op': 'addl'}
    instructions[448] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29, 'op': 'addl'}
    instructions[449] = {5'd3, 4'd6, 4'd0, 16'd867};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29 {'z': 6, 'label': 867, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29, 'op': 'call'}
    instructions[450] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29, 'op': 'addl'}
    instructions[451] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[452] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29, 'op': 'load'}
    instructions[453] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[454] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29, 'op': 'load'}
    instructions[455] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 29, 'op': 'addl'}
    instructions[456] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'store'}
    instructions[457] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'addl'}
    instructions[458] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'store'}
    instructions[459] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'addl'}
    instructions[460] = {5'd0, 4'd8, 4'd0, 16'd41};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'literal': 41, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'literal'}
    instructions[461] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'store'}
    instructions[462] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'addl'}
    instructions[463] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'addl'}
    instructions[464] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'addl'}
    instructions[465] = {5'd3, 4'd6, 4'd0, 16'd479};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'z': 6, 'label': 479, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'call'}
    instructions[466] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'addl'}
    instructions[467] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[468] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'load'}
    instructions[469] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[470] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'load'}
    instructions[471] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 30, 'op': 'addl'}
    instructions[472] = {5'd0, 4'd8, 4'd0, 16'd61568};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 31 {'literal': 61568, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 31, 'op': 'literal'}
    instructions[473] = {5'd6, 4'd8, 4'd8, 16'd762};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 31 {'a': 8, 'literal': 762, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 31, 'op': 'literal_hi'}
    instructions[474] = {5'd10, 4'd0, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 31 {'a': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 31, 'op': 'wait_clocks'}
    instructions[475] = {5'd11, 4'd0, 4'd0, 16'd409};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 26 {'label': 409, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 26, 'op': 'goto'}
    instructions[476] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 9 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 9, 'op': 'addl'}
    instructions[477] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 9 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 9, 'op': 'addl'}
    instructions[478] = {5'd12, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 9 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/temperature.c : 9, 'op': 'return'}
    instructions[479] = {5'd1, 4'd3, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73 {'a': 3, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73, 'op': 'addl'}
    instructions[480] = {5'd2, 4'd0, 4'd3, 16'd6};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'store'}
    instructions[481] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[482] = {5'd2, 4'd0, 4'd3, 16'd7};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'store'}
    instructions[483] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[484] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[485] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[486] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'load'}
    instructions[487] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'store'}
    instructions[488] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[489] = {5'd0, 4'd8, 4'd0, 16'd79};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'literal': 79, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'literal'}
    instructions[490] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[491] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'load'}
    instructions[492] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'store'}
    instructions[493] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[494] = {5'd1, 4'd7, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 4, 'literal': 0, 'z': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[495] = {5'd1, 4'd4, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[496] = {5'd3, 4'd6, 4'd0, 16'd506};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'z': 6, 'label': 506, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'call'}
    instructions[497] = {5'd1, 4'd3, 4'd3, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': -2, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[498] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[499] = {5'd5, 4'd7, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'z': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'load'}
    instructions[500] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[501] = {5'd5, 4'd6, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'z': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'load'}
    instructions[502] = {5'd1, 4'd3, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[503] = {5'd1, 4'd3, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73 {'a': 4, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73, 'op': 'addl'}
    instructions[504] = {5'd1, 4'd4, 4'd7, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73 {'a': 7, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73, 'op': 'addl'}
    instructions[505] = {5'd12, 4'd0, 4'd6, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73 {'a': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73, 'op': 'return'}
    instructions[506] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23, 'op': 'addl'}
    instructions[507] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 24 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 24, 'op': 'literal'}
    instructions[508] = {5'd1, 4'd2, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 24 {'a': 4, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 24, 'op': 'addl'}
    instructions[509] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 24 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 24, 'op': 'store'}
    instructions[510] = {5'd1, 4'd8, 4'd4, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 4, 'literal': -2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'addl'}
    instructions[511] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'addl'}
    instructions[512] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'load'}
    instructions[513] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'store'}
    instructions[514] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'addl'}
    instructions[515] = {5'd1, 4'd8, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 4, 'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'addl'}
    instructions[516] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'addl'}
    instructions[517] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'load'}
    instructions[518] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[519] = {5'd5, 4'd2, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 3, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'load'}
    instructions[520] = {5'd13, 4'd8, 4'd8, 16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 8, 'z': 8, 'b': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'add'}
    instructions[521] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'addl'}
    instructions[522] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'load'}
    instructions[523] = {5'd14, 4'd0, 4'd8, 16'd565};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 29 {'a': 8, 'label': 565, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 29, 'op': 'jmp_if_false'}
    instructions[524] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[525] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[526] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'load'}
    instructions[527] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'store'}
    instructions[528] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[529] = {5'd1, 4'd8, 4'd4, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 4, 'literal': -2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[530] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[531] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'load'}
    instructions[532] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'store'}
    instructions[533] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[534] = {5'd1, 4'd8, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 4, 'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[535] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[536] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'load'}
    instructions[537] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[538] = {5'd5, 4'd2, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'load'}
    instructions[539] = {5'd13, 4'd8, 4'd8, 16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 8, 'z': 8, 'b': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'add'}
    instructions[540] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[541] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'load'}
    instructions[542] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[543] = {5'd5, 4'd0, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'z': 0, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'load'}
    instructions[544] = {5'd15, 4'd0, 4'd0, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 0, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'write'}
    instructions[545] = {5'd1, 4'd3, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[546] = {5'd1, 4'd8, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 4, 'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[547] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[548] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'load'}
    instructions[549] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'store'}
    instructions[550] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[551] = {5'd0, 4'd8, 4'd0, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'literal': 1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'literal'}
    instructions[552] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'store'}
    instructions[553] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[554] = {5'd1, 4'd8, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 4, 'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[555] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[556] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'load'}
    instructions[557] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[558] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'load'}
    instructions[559] = {5'd13, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'add'}
    instructions[560] = {5'd1, 4'd2, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 4, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[561] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'store'}
    instructions[562] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[563] = {5'd5, 4'd8, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'load'}
    instructions[564] = {5'd11, 4'd0, 4'd0, 16'd566};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 29 {'label': 566, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 29, 'op': 'goto'}
    instructions[565] = {5'd11, 4'd0, 4'd0, 16'd567};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 29 {'label': 567, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 29, 'op': 'goto'}
    instructions[566] = {5'd11, 4'd0, 4'd0, 16'd510};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'label': 510, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'goto'}
    instructions[567] = {5'd1, 4'd3, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23 {'a': 4, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23, 'op': 'addl'}
    instructions[568] = {5'd1, 4'd4, 4'd7, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23 {'a': 7, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23, 'op': 'addl'}
    instructions[569] = {5'd12, 4'd0, 4'd6, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23 {'a': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23, 'op': 'return'}
    instructions[570] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 46 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 46, 'op': 'addl'}
    instructions[571] = {5'd1, 4'd8, 4'd4, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 47 {'a': 4, 'literal': -2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 47, 'op': 'addl'}
    instructions[572] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 47 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 47, 'op': 'addl'}
    instructions[573] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 47 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 47, 'op': 'load'}
    instructions[574] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 47 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 47, 'op': 'store'}
    instructions[575] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 47 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 47, 'op': 'addl'}
    instructions[576] = {5'd1, 4'd8, 4'd4, -16'd3};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 47 {'a': 4, 'literal': -3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 47, 'op': 'addl'}
    instructions[577] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 47 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 47, 'op': 'addl'}
    instructions[578] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 47 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 47, 'op': 'load'}
    instructions[579] = {5'd1, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 47 {'a': 8, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 47, 'op': 'addl'}
    instructions[580] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 47 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 47, 'op': 'addl'}
    instructions[581] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 47 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 47, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[582] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 47 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 47, 'op': 'load'}
    instructions[583] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 47 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 47, 'op': 'store'}
    instructions[584] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 48 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 48, 'op': 'addl'}
    instructions[585] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 48 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 48, 'op': 'addl'}
    instructions[586] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 48 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 48, 'op': 'load'}
    instructions[587] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 48 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 48, 'op': 'store'}
    instructions[588] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 48 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 48, 'op': 'addl'}
    instructions[589] = {5'd1, 4'd8, 4'd4, -16'd3};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 48 {'a': 4, 'literal': -3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 48, 'op': 'addl'}
    instructions[590] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 48 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 48, 'op': 'addl'}
    instructions[591] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 48 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 48, 'op': 'load'}
    instructions[592] = {5'd1, 4'd8, 4'd8, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 48 {'a': 8, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 48, 'op': 'addl'}
    instructions[593] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 48 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 48, 'op': 'addl'}
    instructions[594] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 48 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 48, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[595] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 48 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 48, 'op': 'load'}
    instructions[596] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 48 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 48, 'op': 'store'}
    instructions[597] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 46 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 46, 'op': 'addl'}
    instructions[598] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 46 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 46, 'op': 'addl'}
    instructions[599] = {5'd12, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 46 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 46, 'op': 'return'}
    instructions[600] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 9 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 9, 'op': 'addl'}
    instructions[601] = {5'd1, 4'd8, 4'd4, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 10 {'a': 4, 'literal': -2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 10, 'op': 'addl'}
    instructions[602] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 10 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 10, 'op': 'addl'}
    instructions[603] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 10 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 10, 'op': 'load'}
    instructions[604] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 10 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 10, 'op': 'store'}
    instructions[605] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 10 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 10, 'op': 'addl'}
    instructions[606] = {5'd1, 4'd8, 4'd4, -16'd3};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 10 {'a': 4, 'literal': -3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 10, 'op': 'addl'}
    instructions[607] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 10 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 10, 'op': 'addl'}
    instructions[608] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 10 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 10, 'op': 'load'}
    instructions[609] = {5'd1, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 10 {'a': 8, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 10, 'op': 'addl'}
    instructions[610] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 10 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 10, 'op': 'addl'}
    instructions[611] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 10 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 10, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[612] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 10 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 10, 'op': 'load'}
    instructions[613] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 10 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 10, 'op': 'store'}
    instructions[614] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 11 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 11, 'op': 'addl'}
    instructions[615] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 11 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 11, 'op': 'addl'}
    instructions[616] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 11 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 11, 'op': 'load'}
    instructions[617] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 11 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 11, 'op': 'store'}
    instructions[618] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 11 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 11, 'op': 'addl'}
    instructions[619] = {5'd1, 4'd8, 4'd4, -16'd3};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 11 {'a': 4, 'literal': -3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 11, 'op': 'addl'}
    instructions[620] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 11 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 11, 'op': 'addl'}
    instructions[621] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 11 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 11, 'op': 'load'}
    instructions[622] = {5'd1, 4'd8, 4'd8, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 11 {'a': 8, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 11, 'op': 'addl'}
    instructions[623] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 11 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 11, 'op': 'addl'}
    instructions[624] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 11 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 11, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[625] = {5'd5, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 11 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 11, 'op': 'load'}
    instructions[626] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 11 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 11, 'op': 'store'}
    instructions[627] = {5'd0, 4'd8, 4'd0, 16'd61568};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 14 {'literal': 61568, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 14, 'op': 'literal'}
    instructions[628] = {5'd6, 4'd8, 4'd8, 16'd762};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 14 {'a': 8, 'literal': 762, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 14, 'op': 'literal_hi'}
    instructions[629] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 14 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 14, 'op': 'store'}
    instructions[630] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 14 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 14, 'op': 'addl'}
    instructions[631] = {5'd16, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 14 {'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 14, 'op': 'timer_low'}
    instructions[632] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 14 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 14, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[633] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 14 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 14, 'op': 'load'}
    instructions[634] = {5'd17, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 14 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 14, 'op': 'unsigned_greater'}
    instructions[635] = {5'd14, 4'd0, 4'd8, 16'd640};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 14 {'a': 8, 'label': 640, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 14, 'op': 'jmp_if_false'}
    instructions[636] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 14 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 14, 'op': 'addl'}
    instructions[637] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 14 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 14, 'op': 'addl'}
    instructions[638] = {5'd12, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 14 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 14, 'op': 'return'}
    instructions[639] = {5'd11, 4'd0, 4'd0, 16'd640};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 14 {'label': 640, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 14, 'op': 'goto'}
    instructions[640] = {5'd11, 4'd0, 4'd0, 16'd627};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 12 {'label': 627, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 12, 'op': 'goto'}
    instructions[641] = {5'd1, 4'd3, 4'd3, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 19 {'a': 3, 'literal': 2, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 19, 'op': 'addl'}
    instructions[642] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 24 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 24, 'op': 'addl'}
    instructions[643] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 24 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 24, 'op': 'addl'}
    instructions[644] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 24 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 24, 'op': 'load'}
    instructions[645] = {5'd1, 4'd8, 4'd8, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 24 {'a': 8, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 24, 'op': 'addl'}
    instructions[646] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 24 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 24, 'op': 'addl'}
    instructions[647] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 24 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 24, 'op': 'load'}
    instructions[648] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 24 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 24, 'op': 'store'}
    instructions[649] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 24 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 24, 'op': 'addl'}
    instructions[650] = {5'd0, 4'd8, 4'd0, 16'd72};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 24 {'literal': 72, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 24, 'op': 'literal'}
    instructions[651] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 24 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 24, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[652] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 24 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 24, 'op': 'load'}
    instructions[653] = {5'd18, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 24 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 24, 'op': 'or'}
    instructions[654] = {5'd1, 4'd2, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 24 {'a': 4, 'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 24, 'op': 'addl'}
    instructions[655] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 24 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 24, 'op': 'store'}
    instructions[656] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26, 'op': 'store'}
    instructions[657] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26, 'op': 'addl'}
    instructions[658] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26, 'op': 'store'}
    instructions[659] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26, 'op': 'addl'}
    instructions[660] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26, 'op': 'addl'}
    instructions[661] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26, 'op': 'addl'}
    instructions[662] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26, 'op': 'load'}
    instructions[663] = {5'd1, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26 {'a': 8, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26, 'op': 'addl'}
    instructions[664] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26, 'op': 'addl'}
    instructions[665] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26, 'op': 'load'}
    instructions[666] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26, 'op': 'store'}
    instructions[667] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26, 'op': 'addl'}
    instructions[668] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26, 'op': 'literal'}
    instructions[669] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26, 'op': 'store'}
    instructions[670] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26, 'op': 'addl'}
    instructions[671] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26, 'op': 'literal'}
    instructions[672] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26, 'op': 'store'}
    instructions[673] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26, 'op': 'addl'}
    instructions[674] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26, 'op': 'addl'}
    instructions[675] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26, 'op': 'addl'}
    instructions[676] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26, 'op': 'load'}
    instructions[677] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[678] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26, 'op': 'load'}
    instructions[679] = {5'd19, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26, 'op': 'shift_left'}
    instructions[680] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26, 'op': 'store'}
    instructions[681] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26, 'op': 'addl'}
    instructions[682] = {5'd0, 4'd8, 4'd0, 16'd512};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26 {'literal': 512, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26, 'op': 'literal'}
    instructions[683] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[684] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26, 'op': 'load'}
    instructions[685] = {5'd18, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26, 'op': 'or'}
    instructions[686] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[687] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26, 'op': 'load'}
    instructions[688] = {5'd18, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26, 'op': 'or'}
    instructions[689] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26, 'op': 'store'}
    instructions[690] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26, 'op': 'addl'}
    instructions[691] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26, 'op': 'addl'}
    instructions[692] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26, 'op': 'addl'}
    instructions[693] = {5'd3, 4'd6, 4'd0, 16'd788};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26 {'z': 6, 'label': 788, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26, 'op': 'call'}
    instructions[694] = {5'd1, 4'd3, 4'd3, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26 {'a': 3, 'literal': -2, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26, 'op': 'addl'}
    instructions[695] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[696] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26, 'op': 'load'}
    instructions[697] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[698] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26, 'op': 'load'}
    instructions[699] = {5'd0, 4'd2, 4'd0, 16'd106};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26 {'literal': 106, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26, 'op': 'literal'}
    instructions[700] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 26, 'op': 'load'}
    instructions[701] = {5'd0, 4'd8, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27 {'literal': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27, 'op': 'literal'}
    instructions[702] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27, 'op': 'store'}
    instructions[703] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27, 'op': 'addl'}
    instructions[704] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27, 'op': 'store'}
    instructions[705] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27, 'op': 'addl'}
    instructions[706] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27, 'op': 'store'}
    instructions[707] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27, 'op': 'addl'}
    instructions[708] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27, 'op': 'addl'}
    instructions[709] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27, 'op': 'addl'}
    instructions[710] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27, 'op': 'load'}
    instructions[711] = {5'd1, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27 {'a': 8, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27, 'op': 'addl'}
    instructions[712] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27, 'op': 'addl'}
    instructions[713] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27, 'op': 'load'}
    instructions[714] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27, 'op': 'store'}
    instructions[715] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27, 'op': 'addl'}
    instructions[716] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27, 'op': 'literal'}
    instructions[717] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27, 'op': 'store'}
    instructions[718] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27, 'op': 'addl'}
    instructions[719] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27, 'op': 'addl'}
    instructions[720] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27, 'op': 'addl'}
    instructions[721] = {5'd3, 4'd6, 4'd0, 16'd822};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27 {'z': 6, 'label': 822, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27, 'op': 'call'}
    instructions[722] = {5'd1, 4'd3, 4'd3, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27 {'a': 3, 'literal': -2, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27, 'op': 'addl'}
    instructions[723] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[724] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27, 'op': 'load'}
    instructions[725] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[726] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27, 'op': 'load'}
    instructions[727] = {5'd0, 4'd2, 4'd0, 16'd39};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27 {'literal': 39, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27, 'op': 'literal'}
    instructions[728] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27, 'op': 'load'}
    instructions[729] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[730] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27, 'op': 'load'}
    instructions[731] = {5'd19, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27, 'op': 'shift_left'}
    instructions[732] = {5'd1, 4'd2, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27, 'op': 'addl'}
    instructions[733] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 27, 'op': 'store'}
    instructions[734] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28, 'op': 'store'}
    instructions[735] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28, 'op': 'addl'}
    instructions[736] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28, 'op': 'store'}
    instructions[737] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28, 'op': 'addl'}
    instructions[738] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28, 'op': 'addl'}
    instructions[739] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28, 'op': 'addl'}
    instructions[740] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28, 'op': 'load'}
    instructions[741] = {5'd1, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28 {'a': 8, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28, 'op': 'addl'}
    instructions[742] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28, 'op': 'addl'}
    instructions[743] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28, 'op': 'load'}
    instructions[744] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28, 'op': 'store'}
    instructions[745] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28, 'op': 'addl'}
    instructions[746] = {5'd0, 4'd8, 4'd0, 16'd3072};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28 {'literal': 3072, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28, 'op': 'literal'}
    instructions[747] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28, 'op': 'store'}
    instructions[748] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28, 'op': 'addl'}
    instructions[749] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28, 'op': 'addl'}
    instructions[750] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28, 'op': 'addl'}
    instructions[751] = {5'd3, 4'd6, 4'd0, 16'd822};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28 {'z': 6, 'label': 822, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28, 'op': 'call'}
    instructions[752] = {5'd1, 4'd3, 4'd3, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28 {'a': 3, 'literal': -2, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28, 'op': 'addl'}
    instructions[753] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[754] = {5'd5, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28, 'op': 'load'}
    instructions[755] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[756] = {5'd5, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28, 'op': 'load'}
    instructions[757] = {5'd0, 4'd2, 4'd0, 16'd39};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28 {'literal': 39, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28, 'op': 'literal'}
    instructions[758] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28, 'op': 'load'}
    instructions[759] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28, 'op': 'store'}
    instructions[760] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28, 'op': 'addl'}
    instructions[761] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28, 'op': 'addl'}
    instructions[762] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28, 'op': 'addl'}
    instructions[763] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28, 'op': 'load'}
    instructions[764] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[765] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28, 'op': 'load'}
    instructions[766] = {5'd18, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28, 'op': 'or'}
    instructions[767] = {5'd1, 4'd2, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28, 'op': 'addl'}
    instructions[768] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 28, 'op': 'store'}
    instructions[769] = {5'd0, 4'd8, 4'd0, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 29 {'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 29, 'op': 'literal'}
    instructions[770] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 29 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 29, 'op': 'store'}
    instructions[771] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 29 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 29, 'op': 'addl'}
    instructions[772] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 29 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 29, 'op': 'addl'}
    instructions[773] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 29 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 29, 'op': 'addl'}
    instructions[774] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 29 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 29, 'op': 'load'}
    instructions[775] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 29 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 29, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[776] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 29 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 29, 'op': 'load'}
    instructions[777] = {5'd20, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 29 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 29, 'op': 'unsigned_shift_right'}
    instructions[778] = {5'd1, 4'd2, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 29 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 29, 'op': 'addl'}
    instructions[779] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 29 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 29, 'op': 'store'}
    instructions[780] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 30 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 30, 'op': 'addl'}
    instructions[781] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 30 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 30, 'op': 'addl'}
    instructions[782] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 30 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 30, 'op': 'load'}
    instructions[783] = {5'd0, 4'd2, 4'd0, 16'd37};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 30 {'literal': 37, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 30, 'op': 'literal'}
    instructions[784] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 30 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 30, 'op': 'store'}
    instructions[785] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 30 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 30, 'op': 'addl'}
    instructions[786] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 30 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 30, 'op': 'addl'}
    instructions[787] = {5'd12, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 30 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/adt7420.h : 30, 'op': 'return'}
    instructions[788] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 52 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 52, 'op': 'addl'}
    instructions[789] = {5'd1, 4'd8, 4'd4, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 57 {'a': 4, 'literal': -2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 57, 'op': 'addl'}
    instructions[790] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 57 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 57, 'op': 'addl'}
    instructions[791] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 57 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 57, 'op': 'load'}
    instructions[792] = {5'd1, 4'd8, 4'd8, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 57 {'a': 8, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 57, 'op': 'addl'}
    instructions[793] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 57 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 57, 'op': 'addl'}
    instructions[794] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 57 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 57, 'op': 'load'}
    instructions[795] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 57 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 57, 'op': 'store'}
    instructions[796] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 57 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 57, 'op': 'addl'}
    instructions[797] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 57 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 57, 'op': 'addl'}
    instructions[798] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 57 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 57, 'op': 'addl'}
    instructions[799] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 57 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 57, 'op': 'load'}
    instructions[800] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 57 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 57, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[801] = {5'd5, 4'd0, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 57 {'a': 3, 'z': 0, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 57, 'op': 'load'}
    instructions[802] = {5'd15, 4'd0, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 57 {'a': 0, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 57, 'op': 'write'}
    instructions[803] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 57 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 57, 'op': 'addl'}
    instructions[804] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 58 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 58, 'op': 'literal'}
    instructions[805] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 58 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 58, 'op': 'store'}
    instructions[806] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 58 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 58, 'op': 'addl'}
    instructions[807] = {5'd1, 4'd8, 4'd4, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 58 {'a': 4, 'literal': -2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 58, 'op': 'addl'}
    instructions[808] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 58 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 58, 'op': 'addl'}
    instructions[809] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 58 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 58, 'op': 'load'}
    instructions[810] = {5'd1, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 58 {'a': 8, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 58, 'op': 'addl'}
    instructions[811] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 58 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 58, 'op': 'addl'}
    instructions[812] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 58 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 58, 'op': 'load'}
    instructions[813] = {5'd21, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 58 {'a': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 58, 'op': 'read'}
    instructions[814] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 58 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 58, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[815] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 58 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 58, 'op': 'load'}
    instructions[816] = {5'd22, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 58 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 58, 'op': 'and'}
    instructions[817] = {5'd0, 4'd2, 4'd0, 16'd106};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 58 {'literal': 106, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 58, 'op': 'literal'}
    instructions[818] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 58 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 58, 'op': 'store'}
    instructions[819] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 58 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 58, 'op': 'addl'}
    instructions[820] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 58 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 58, 'op': 'addl'}
    instructions[821] = {5'd12, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 58 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 58, 'op': 'return'}
    instructions[822] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 62 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 62, 'op': 'addl'}
    instructions[823] = {5'd0, 4'd8, 4'd0, 16'd256};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 66 {'literal': 256, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 66, 'op': 'literal'}
    instructions[824] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 66 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 66, 'op': 'store'}
    instructions[825] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 66 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 66, 'op': 'addl'}
    instructions[826] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 66 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 66, 'op': 'addl'}
    instructions[827] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 66 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 66, 'op': 'addl'}
    instructions[828] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 66 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 66, 'op': 'load'}
    instructions[829] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 66 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 66, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[830] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 66 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 66, 'op': 'load'}
    instructions[831] = {5'd18, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 66 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 66, 'op': 'or'}
    instructions[832] = {5'd1, 4'd2, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 66 {'a': 4, 'literal': -1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 66, 'op': 'addl'}
    instructions[833] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 66 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 66, 'op': 'store'}
    instructions[834] = {5'd1, 4'd8, 4'd4, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 67 {'a': 4, 'literal': -2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 67, 'op': 'addl'}
    instructions[835] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 67 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 67, 'op': 'addl'}
    instructions[836] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 67 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 67, 'op': 'load'}
    instructions[837] = {5'd1, 4'd8, 4'd8, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 67 {'a': 8, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 67, 'op': 'addl'}
    instructions[838] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 67 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 67, 'op': 'addl'}
    instructions[839] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 67 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 67, 'op': 'load'}
    instructions[840] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 67 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 67, 'op': 'store'}
    instructions[841] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 67 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 67, 'op': 'addl'}
    instructions[842] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 67 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 67, 'op': 'addl'}
    instructions[843] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 67 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 67, 'op': 'addl'}
    instructions[844] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 67 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 67, 'op': 'load'}
    instructions[845] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 67 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 67, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[846] = {5'd5, 4'd0, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 67 {'a': 3, 'z': 0, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 67, 'op': 'load'}
    instructions[847] = {5'd15, 4'd0, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 67 {'a': 0, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 67, 'op': 'write'}
    instructions[848] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 67 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 67, 'op': 'addl'}
    instructions[849] = {5'd0, 4'd8, 4'd0, 16'd255};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 68 {'literal': 255, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 68, 'op': 'literal'}
    instructions[850] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 68 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 68, 'op': 'store'}
    instructions[851] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 68 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 68, 'op': 'addl'}
    instructions[852] = {5'd1, 4'd8, 4'd4, -16'd2};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 68 {'a': 4, 'literal': -2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 68, 'op': 'addl'}
    instructions[853] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 68 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 68, 'op': 'addl'}
    instructions[854] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 68 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 68, 'op': 'load'}
    instructions[855] = {5'd1, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 68 {'a': 8, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 68, 'op': 'addl'}
    instructions[856] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 68 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 68, 'op': 'addl'}
    instructions[857] = {5'd5, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 68 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 68, 'op': 'load'}
    instructions[858] = {5'd21, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 68 {'a': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 68, 'op': 'read'}
    instructions[859] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 68 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 68, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[860] = {5'd5, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 68 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 68, 'op': 'load'}
    instructions[861] = {5'd22, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 68 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 68, 'op': 'and'}
    instructions[862] = {5'd0, 4'd2, 4'd0, 16'd39};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 68 {'literal': 39, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 68, 'op': 'literal'}
    instructions[863] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 68 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 68, 'op': 'store'}
    instructions[864] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 68 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 68, 'op': 'addl'}
    instructions[865] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 68 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 68, 'op': 'addl'}
    instructions[866] = {5'd12, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 68 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/temperature/i2c.h : 68, 'op': 'return'}
    instructions[867] = {5'd1, 4'd3, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 165 {'a': 3, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 165, 'op': 'addl'}
    instructions[868] = {5'd2, 4'd0, 4'd3, 16'd6};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 166 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 166, 'op': 'store'}
    instructions[869] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 166 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 166, 'op': 'addl'}
    instructions[870] = {5'd2, 4'd0, 4'd3, 16'd7};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 166 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 166, 'op': 'store'}
    instructions[871] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 166 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 166, 'op': 'addl'}
    instructions[872] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 166 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 166, 'op': 'addl'}
    instructions[873] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 166 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 166, 'op': 'addl'}
    instructions[874] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 166 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 166, 'op': 'load'}
    instructions[875] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 166 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 166, 'op': 'store'}
    instructions[876] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 166 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 166, 'op': 'addl'}
    instructions[877] = {5'd0, 4'd8, 4'd0, 16'd79};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 166 {'literal': 79, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 166, 'op': 'literal'}
    instructions[878] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 166 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 166, 'op': 'addl'}
    instructions[879] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 166 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 166, 'op': 'load'}
    instructions[880] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 166 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 166, 'op': 'store'}
    instructions[881] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 166 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 166, 'op': 'addl'}
    instructions[882] = {5'd1, 4'd7, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 166 {'a': 4, 'literal': 0, 'z': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 166, 'op': 'addl'}
    instructions[883] = {5'd1, 4'd4, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 166 {'a': 3, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 166, 'op': 'addl'}
    instructions[884] = {5'd3, 4'd6, 4'd0, 16'd894};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 166 {'z': 6, 'label': 894, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 166, 'op': 'call'}
    instructions[885] = {5'd1, 4'd3, 4'd3, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 166 {'a': 3, 'literal': -2, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 166, 'op': 'addl'}
    instructions[886] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 166 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 166, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[887] = {5'd5, 4'd7, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 166 {'a': 3, 'z': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 166, 'op': 'load'}
    instructions[888] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 166 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 166, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[889] = {5'd5, 4'd6, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 166 {'a': 3, 'z': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 166, 'op': 'load'}
    instructions[890] = {5'd1, 4'd3, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 166 {'a': 3, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 166, 'op': 'addl'}
    instructions[891] = {5'd1, 4'd3, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 165 {'a': 4, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 165, 'op': 'addl'}
    instructions[892] = {5'd1, 4'd4, 4'd7, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 165 {'a': 7, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 165, 'op': 'addl'}
    instructions[893] = {5'd12, 4'd0, 4'd6, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 165 {'a': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 165, 'op': 'return'}
    instructions[894] = {5'd1, 4'd3, 4'd3, 16'd3};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 79 {'a': 3, 'literal': 3, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 79, 'op': 'addl'}
    instructions[895] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 81 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 81, 'op': 'literal'}
    instructions[896] = {5'd1, 4'd2, 4'd4, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 81 {'a': 4, 'literal': 1, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 81, 'op': 'addl'}
    instructions[897] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 81 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 81, 'op': 'store'}
    instructions[898] = {5'd0, 4'd8, 4'd0, 16'd48160};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 82 {'literal': 48160, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 82, 'op': 'literal'}
    instructions[899] = {5'd6, 4'd8, 4'd8, 16'd19646};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 82 {'a': 8, 'literal': 19646, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 82, 'op': 'literal_hi'}
    instructions[900] = {5'd1, 4'd2, 4'd4, 16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 82 {'a': 4, 'literal': 2, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 82, 'op': 'addl'}
    instructions[901] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 82 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 82, 'op': 'store'}
    instructions[902] = {5'd2, 4'd0, 4'd3, 16'd6};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84, 'op': 'store'}
    instructions[903] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84, 'op': 'addl'}
    instructions[904] = {5'd2, 4'd0, 4'd3, 16'd7};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84, 'op': 'store'}
    instructions[905] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84, 'op': 'addl'}
    instructions[906] = {5'd1, 4'd8, 4'd4, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84 {'a': 4, 'literal': -2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84, 'op': 'addl'}
    instructions[907] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84, 'op': 'addl'}
    instructions[908] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84, 'op': 'load'}
    instructions[909] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84, 'op': 'store'}
    instructions[910] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84, 'op': 'addl'}
    instructions[911] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84, 'op': 'literal'}
    instructions[912] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84, 'op': 'store'}
    instructions[913] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84, 'op': 'addl'}
    instructions[914] = {5'd1, 4'd7, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84 {'a': 4, 'literal': 0, 'z': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84, 'op': 'addl'}
    instructions[915] = {5'd1, 4'd4, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84 {'a': 3, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84, 'op': 'addl'}
    instructions[916] = {5'd3, 4'd6, 4'd0, 16'd1225};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84 {'z': 6, 'label': 1225, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84, 'op': 'call'}
    instructions[917] = {5'd1, 4'd3, 4'd3, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84 {'a': 3, 'literal': -2, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84, 'op': 'addl'}
    instructions[918] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[919] = {5'd5, 4'd7, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84 {'a': 3, 'z': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84, 'op': 'load'}
    instructions[920] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[921] = {5'd5, 4'd6, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84 {'a': 3, 'z': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84, 'op': 'load'}
    instructions[922] = {5'd0, 4'd2, 4'd0, 16'd80};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84 {'literal': 80, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84, 'op': 'literal'}
    instructions[923] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84, 'op': 'load'}
    instructions[924] = {5'd14, 4'd0, 4'd8, 16'd947};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84 {'a': 8, 'label': 947, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84, 'op': 'jmp_if_false'}
    instructions[925] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 85 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 85, 'op': 'addl'}
    instructions[926] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 85 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 85, 'op': 'addl'}
    instructions[927] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 85 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 85, 'op': 'load'}
    instructions[928] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 85 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 85, 'op': 'store'}
    instructions[929] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 85 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 85, 'op': 'addl'}
    instructions[930] = {5'd0, 4'd8, 4'd0, 16'd45};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 85 {'literal': 45, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 85, 'op': 'literal'}
    instructions[931] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 85 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 85, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[932] = {5'd5, 4'd0, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 85 {'a': 3, 'z': 0, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 85, 'op': 'load'}
    instructions[933] = {5'd15, 4'd0, 4'd0, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 85 {'a': 0, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 85, 'op': 'write'}
    instructions[934] = {5'd1, 4'd3, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 85 {'a': 3, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 85, 'op': 'addl'}
    instructions[935] = {5'd1, 4'd8, 4'd4, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 86 {'a': 4, 'literal': -2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 86, 'op': 'addl'}
    instructions[936] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 86 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 86, 'op': 'addl'}
    instructions[937] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 86 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 86, 'op': 'load'}
    instructions[938] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 86 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 86, 'op': 'store'}
    instructions[939] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 86 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 86, 'op': 'addl'}
    instructions[940] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 86 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 86, 'op': 'literal'}
    instructions[941] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 86 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 86, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[942] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 86 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 86, 'op': 'load'}
    instructions[943] = {5'd23, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 86 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 86, 'op': 'float_subtract'}
    instructions[944] = {5'd1, 4'd2, 4'd4, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 86 {'a': 4, 'literal': -2, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 86, 'op': 'addl'}
    instructions[945] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 86 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 86, 'op': 'store'}
    instructions[946] = {5'd11, 4'd0, 4'd0, 16'd947};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84 {'label': 947, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 84, 'op': 'goto'}
    instructions[947] = {5'd2, 4'd0, 4'd3, 16'd6};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89, 'op': 'store'}
    instructions[948] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89, 'op': 'addl'}
    instructions[949] = {5'd2, 4'd0, 4'd3, 16'd7};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89, 'op': 'store'}
    instructions[950] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89, 'op': 'addl'}
    instructions[951] = {5'd1, 4'd8, 4'd4, 16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89 {'a': 4, 'literal': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89, 'op': 'addl'}
    instructions[952] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89, 'op': 'addl'}
    instructions[953] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89, 'op': 'load'}
    instructions[954] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89, 'op': 'store'}
    instructions[955] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89, 'op': 'addl'}
    instructions[956] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89, 'op': 'literal'}
    instructions[957] = {5'd6, 4'd8, 4'd8, 16'd16256};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89 {'a': 8, 'literal': 16256, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89, 'op': 'literal_hi'}
    instructions[958] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89, 'op': 'store'}
    instructions[959] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89, 'op': 'addl'}
    instructions[960] = {5'd1, 4'd7, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89 {'a': 4, 'literal': 0, 'z': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89, 'op': 'addl'}
    instructions[961] = {5'd1, 4'd4, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89 {'a': 3, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89, 'op': 'addl'}
    instructions[962] = {5'd3, 4'd6, 4'd0, 16'd1288};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89 {'z': 6, 'label': 1288, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89, 'op': 'call'}
    instructions[963] = {5'd1, 4'd3, 4'd3, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89 {'a': 3, 'literal': -2, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89, 'op': 'addl'}
    instructions[964] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[965] = {5'd5, 4'd7, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89 {'a': 3, 'z': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89, 'op': 'load'}
    instructions[966] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[967] = {5'd5, 4'd6, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89 {'a': 3, 'z': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89, 'op': 'load'}
    instructions[968] = {5'd0, 4'd2, 4'd0, 16'd105};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89 {'literal': 105, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89, 'op': 'literal'}
    instructions[969] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89, 'op': 'load'}
    instructions[970] = {5'd14, 4'd0, 4'd8, 16'd1088};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 103 {'a': 8, 'label': 1088, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 103, 'op': 'jmp_if_false'}
    instructions[971] = {5'd1, 4'd8, 4'd4, 16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 90 {'a': 4, 'literal': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 90, 'op': 'addl'}
    instructions[972] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 90 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 90, 'op': 'addl'}
    instructions[973] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 90 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 90, 'op': 'load'}
    instructions[974] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 90 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 90, 'op': 'store'}
    instructions[975] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 90 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 90, 'op': 'addl'}
    instructions[976] = {5'd1, 4'd8, 4'd4, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 90 {'a': 4, 'literal': -2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 90, 'op': 'addl'}
    instructions[977] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 90 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 90, 'op': 'addl'}
    instructions[978] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 90 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 90, 'op': 'load'}
    instructions[979] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 90 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 90, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[980] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 90 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 90, 'op': 'load'}
    instructions[981] = {5'd24, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 90 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 90, 'op': 'float_divide'}
    instructions[982] = {5'd7, 4'd8, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 90 {'a': 8, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 90, 'op': 'a_lo'}
    instructions[983] = {5'd25, 4'd0, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 90 {'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 90, 'op': 'float_to_int'}
    instructions[984] = {5'd7, 4'd8, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 90 {'a': 8, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 90, 'op': 'a_lo'}
    instructions[985] = {5'd1, 4'd2, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 90 {'a': 4, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 90, 'op': 'addl'}
    instructions[986] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 90 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 90, 'op': 'store'}
    instructions[987] = {5'd2, 4'd0, 4'd3, 16'd6};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91, 'op': 'store'}
    instructions[988] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91, 'op': 'addl'}
    instructions[989] = {5'd2, 4'd0, 4'd3, 16'd7};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91, 'op': 'store'}
    instructions[990] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91, 'op': 'addl'}
    instructions[991] = {5'd1, 4'd8, 4'd4, 16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91 {'a': 4, 'literal': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91, 'op': 'addl'}
    instructions[992] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91, 'op': 'addl'}
    instructions[993] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91, 'op': 'load'}
    instructions[994] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91, 'op': 'store'}
    instructions[995] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91, 'op': 'addl'}
    instructions[996] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91, 'op': 'literal'}
    instructions[997] = {5'd6, 4'd8, 4'd8, 16'd16672};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91 {'a': 8, 'literal': 16672, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91, 'op': 'literal_hi'}
    instructions[998] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91, 'op': 'store'}
    instructions[999] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91, 'op': 'addl'}
    instructions[1000] = {5'd1, 4'd7, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91 {'a': 4, 'literal': 0, 'z': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91, 'op': 'addl'}
    instructions[1001] = {5'd1, 4'd4, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91 {'a': 3, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91, 'op': 'addl'}
    instructions[1002] = {5'd3, 4'd6, 4'd0, 16'd1225};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91 {'z': 6, 'label': 1225, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91, 'op': 'call'}
    instructions[1003] = {5'd1, 4'd3, 4'd3, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91 {'a': 3, 'literal': -2, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91, 'op': 'addl'}
    instructions[1004] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1005] = {5'd5, 4'd7, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91 {'a': 3, 'z': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91, 'op': 'load'}
    instructions[1006] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1007] = {5'd5, 4'd6, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91 {'a': 3, 'z': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91, 'op': 'load'}
    instructions[1008] = {5'd0, 4'd2, 4'd0, 16'd80};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91 {'literal': 80, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91, 'op': 'literal'}
    instructions[1009] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91, 'op': 'load'}
    instructions[1010] = {5'd14, 4'd0, 4'd8, 16'd1015};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91 {'a': 8, 'label': 1015, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91, 'op': 'jmp_if_false'}
    instructions[1011] = {5'd0, 4'd8, 4'd0, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 92 {'literal': 1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 92, 'op': 'literal'}
    instructions[1012] = {5'd1, 4'd2, 4'd4, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 92 {'a': 4, 'literal': 1, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 92, 'op': 'addl'}
    instructions[1013] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 92 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 92, 'op': 'store'}
    instructions[1014] = {5'd11, 4'd0, 4'd0, 16'd1028};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91 {'label': 1028, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 91, 'op': 'goto'}
    instructions[1015] = {5'd1, 4'd8, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 94 {'a': 4, 'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 94, 'op': 'addl'}
    instructions[1016] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 94 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 94, 'op': 'addl'}
    instructions[1017] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 94 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 94, 'op': 'load'}
    instructions[1018] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 94 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 94, 'op': 'store'}
    instructions[1019] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 94 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 94, 'op': 'addl'}
    instructions[1020] = {5'd1, 4'd8, 4'd4, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 94 {'a': 4, 'literal': 1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 94, 'op': 'addl'}
    instructions[1021] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 94 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 94, 'op': 'addl'}
    instructions[1022] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 94 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 94, 'op': 'load'}
    instructions[1023] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 94 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 94, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1024] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 94 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 94, 'op': 'load'}
    instructions[1025] = {5'd18, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 94 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 94, 'op': 'or'}
    instructions[1026] = {5'd1, 4'd2, 4'd4, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 94 {'a': 4, 'literal': 1, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 94, 'op': 'addl'}
    instructions[1027] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 94 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 94, 'op': 'store'}
    instructions[1028] = {5'd1, 4'd8, 4'd4, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 96 {'a': 4, 'literal': 1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 96, 'op': 'addl'}
    instructions[1029] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 96 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 96, 'op': 'addl'}
    instructions[1030] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 96 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 96, 'op': 'load'}
    instructions[1031] = {5'd14, 4'd0, 4'd8, 16'd1051};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 96 {'a': 8, 'label': 1051, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 96, 'op': 'jmp_if_false'}
    instructions[1032] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 97 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 97, 'op': 'addl'}
    instructions[1033] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 97 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 97, 'op': 'addl'}
    instructions[1034] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 97 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 97, 'op': 'load'}
    instructions[1035] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 97 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 97, 'op': 'store'}
    instructions[1036] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 97 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 97, 'op': 'addl'}
    instructions[1037] = {5'd0, 4'd8, 4'd0, 16'd48};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 97 {'literal': 48, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 97, 'op': 'literal'}
    instructions[1038] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 97 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 97, 'op': 'store'}
    instructions[1039] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 97 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 97, 'op': 'addl'}
    instructions[1040] = {5'd1, 4'd8, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 97 {'a': 4, 'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 97, 'op': 'addl'}
    instructions[1041] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 97 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 97, 'op': 'addl'}
    instructions[1042] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 97 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 97, 'op': 'load'}
    instructions[1043] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 97 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 97, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1044] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 97 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 97, 'op': 'load'}
    instructions[1045] = {5'd13, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 97 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 97, 'op': 'add'}
    instructions[1046] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 97 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 97, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1047] = {5'd5, 4'd0, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 97 {'a': 3, 'z': 0, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 97, 'op': 'load'}
    instructions[1048] = {5'd15, 4'd0, 4'd0, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 97 {'a': 0, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 97, 'op': 'write'}
    instructions[1049] = {5'd1, 4'd3, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 97 {'a': 3, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 97, 'op': 'addl'}
    instructions[1050] = {5'd11, 4'd0, 4'd0, 16'd1051};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 96 {'label': 1051, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 96, 'op': 'goto'}
    instructions[1051] = {5'd1, 4'd8, 4'd4, 16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99 {'a': 4, 'literal': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99, 'op': 'addl'}
    instructions[1052] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99, 'op': 'addl'}
    instructions[1053] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99, 'op': 'load'}
    instructions[1054] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99, 'op': 'store'}
    instructions[1055] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99, 'op': 'addl'}
    instructions[1056] = {5'd1, 4'd8, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99 {'a': 4, 'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99, 'op': 'addl'}
    instructions[1057] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99, 'op': 'addl'}
    instructions[1058] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99, 'op': 'load'}
    instructions[1059] = {5'd7, 4'd8, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99 {'a': 8, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99, 'op': 'a_lo'}
    instructions[1060] = {5'd8, 4'd0, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99 {'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99, 'op': 'int_to_float'}
    instructions[1061] = {5'd7, 4'd8, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99 {'a': 8, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99, 'op': 'a_lo'}
    instructions[1062] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1063] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99, 'op': 'load'}
    instructions[1064] = {5'd9, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99, 'op': 'float_multiply'}
    instructions[1065] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99, 'op': 'store'}
    instructions[1066] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99, 'op': 'addl'}
    instructions[1067] = {5'd1, 4'd8, 4'd4, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99 {'a': 4, 'literal': -2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99, 'op': 'addl'}
    instructions[1068] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99, 'op': 'addl'}
    instructions[1069] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99, 'op': 'load'}
    instructions[1070] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1071] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99, 'op': 'load'}
    instructions[1072] = {5'd23, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99, 'op': 'float_subtract'}
    instructions[1073] = {5'd1, 4'd2, 4'd4, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99 {'a': 4, 'literal': -2, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99, 'op': 'addl'}
    instructions[1074] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 99, 'op': 'store'}
    instructions[1075] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 100 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 100, 'op': 'literal'}
    instructions[1076] = {5'd6, 4'd8, 4'd8, 16'd16672};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 100 {'a': 8, 'literal': 16672, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 100, 'op': 'literal_hi'}
    instructions[1077] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 100 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 100, 'op': 'store'}
    instructions[1078] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 100 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 100, 'op': 'addl'}
    instructions[1079] = {5'd1, 4'd8, 4'd4, 16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 100 {'a': 4, 'literal': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 100, 'op': 'addl'}
    instructions[1080] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 100 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 100, 'op': 'addl'}
    instructions[1081] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 100 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 100, 'op': 'load'}
    instructions[1082] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 100 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 100, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1083] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 100 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 100, 'op': 'load'}
    instructions[1084] = {5'd24, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 100 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 100, 'op': 'float_divide'}
    instructions[1085] = {5'd1, 4'd2, 4'd4, 16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 100 {'a': 4, 'literal': 2, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 100, 'op': 'addl'}
    instructions[1086] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 100 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 100, 'op': 'store'}
    instructions[1087] = {5'd11, 4'd0, 4'd0, 16'd1089};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 103 {'label': 1089, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 103, 'op': 'goto'}
    instructions[1088] = {5'd11, 4'd0, 4'd0, 16'd1090};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 103 {'label': 1090, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 103, 'op': 'goto'}
    instructions[1089] = {5'd11, 4'd0, 4'd0, 16'd947};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89 {'label': 947, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 89, 'op': 'goto'}
    instructions[1090] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 103 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 103, 'op': 'addl'}
    instructions[1091] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 103 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 103, 'op': 'addl'}
    instructions[1092] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 103 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 103, 'op': 'load'}
    instructions[1093] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 103 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 103, 'op': 'store'}
    instructions[1094] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 103 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 103, 'op': 'addl'}
    instructions[1095] = {5'd0, 4'd8, 4'd0, 16'd46};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 103 {'literal': 46, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 103, 'op': 'literal'}
    instructions[1096] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 103 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 103, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1097] = {5'd5, 4'd0, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 103 {'a': 3, 'z': 0, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 103, 'op': 'load'}
    instructions[1098] = {5'd15, 4'd0, 4'd0, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 103 {'a': 0, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 103, 'op': 'write'}
    instructions[1099] = {5'd1, 4'd3, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 103 {'a': 3, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 103, 'op': 'addl'}
    instructions[1100] = {5'd2, 4'd0, 4'd3, 16'd6};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105, 'op': 'store'}
    instructions[1101] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105, 'op': 'addl'}
    instructions[1102] = {5'd2, 4'd0, 4'd3, 16'd7};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105, 'op': 'store'}
    instructions[1103] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105, 'op': 'addl'}
    instructions[1104] = {5'd1, 4'd8, 4'd4, 16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105 {'a': 4, 'literal': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105, 'op': 'addl'}
    instructions[1105] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105, 'op': 'addl'}
    instructions[1106] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105, 'op': 'load'}
    instructions[1107] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105, 'op': 'store'}
    instructions[1108] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105, 'op': 'addl'}
    instructions[1109] = {5'd0, 4'd8, 4'd0, 16'd52343};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105 {'literal': 52343, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105, 'op': 'literal'}
    instructions[1110] = {5'd6, 4'd8, 4'd8, 16'd12843};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105 {'a': 8, 'literal': 12843, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105, 'op': 'literal_hi'}
    instructions[1111] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105, 'op': 'store'}
    instructions[1112] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105, 'op': 'addl'}
    instructions[1113] = {5'd1, 4'd7, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105 {'a': 4, 'literal': 0, 'z': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105, 'op': 'addl'}
    instructions[1114] = {5'd1, 4'd4, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105 {'a': 3, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105, 'op': 'addl'}
    instructions[1115] = {5'd3, 4'd6, 4'd0, 16'd1351};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105 {'z': 6, 'label': 1351, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105, 'op': 'call'}
    instructions[1116] = {5'd1, 4'd3, 4'd3, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105 {'a': 3, 'literal': -2, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105, 'op': 'addl'}
    instructions[1117] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1118] = {5'd5, 4'd7, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105 {'a': 3, 'z': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105, 'op': 'load'}
    instructions[1119] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1120] = {5'd5, 4'd6, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105 {'a': 3, 'z': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105, 'op': 'load'}
    instructions[1121] = {5'd0, 4'd2, 4'd0, 16'd82};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105 {'literal': 82, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105, 'op': 'literal'}
    instructions[1122] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105, 'op': 'load'}
    instructions[1123] = {5'd14, 4'd0, 4'd8, 16'd1220};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 112 {'a': 8, 'label': 1220, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 112, 'op': 'jmp_if_false'}
    instructions[1124] = {5'd1, 4'd8, 4'd4, 16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 106 {'a': 4, 'literal': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 106, 'op': 'addl'}
    instructions[1125] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 106 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 106, 'op': 'addl'}
    instructions[1126] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 106 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 106, 'op': 'load'}
    instructions[1127] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 106 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 106, 'op': 'store'}
    instructions[1128] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 106 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 106, 'op': 'addl'}
    instructions[1129] = {5'd1, 4'd8, 4'd4, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 106 {'a': 4, 'literal': -2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 106, 'op': 'addl'}
    instructions[1130] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 106 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 106, 'op': 'addl'}
    instructions[1131] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 106 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 106, 'op': 'load'}
    instructions[1132] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 106 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 106, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1133] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 106 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 106, 'op': 'load'}
    instructions[1134] = {5'd24, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 106 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 106, 'op': 'float_divide'}
    instructions[1135] = {5'd7, 4'd8, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 106 {'a': 8, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 106, 'op': 'a_lo'}
    instructions[1136] = {5'd25, 4'd0, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 106 {'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 106, 'op': 'float_to_int'}
    instructions[1137] = {5'd7, 4'd8, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 106 {'a': 8, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 106, 'op': 'a_lo'}
    instructions[1138] = {5'd1, 4'd2, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 106 {'a': 4, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 106, 'op': 'addl'}
    instructions[1139] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 106 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 106, 'op': 'store'}
    instructions[1140] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 107 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 107, 'op': 'addl'}
    instructions[1141] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 107 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 107, 'op': 'addl'}
    instructions[1142] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 107 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 107, 'op': 'load'}
    instructions[1143] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 107 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 107, 'op': 'store'}
    instructions[1144] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 107 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 107, 'op': 'addl'}
    instructions[1145] = {5'd0, 4'd8, 4'd0, 16'd48};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 107 {'literal': 48, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 107, 'op': 'literal'}
    instructions[1146] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 107 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 107, 'op': 'store'}
    instructions[1147] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 107 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 107, 'op': 'addl'}
    instructions[1148] = {5'd1, 4'd8, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 107 {'a': 4, 'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 107, 'op': 'addl'}
    instructions[1149] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 107 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 107, 'op': 'addl'}
    instructions[1150] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 107 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 107, 'op': 'load'}
    instructions[1151] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 107 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 107, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1152] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 107 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 107, 'op': 'load'}
    instructions[1153] = {5'd13, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 107 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 107, 'op': 'add'}
    instructions[1154] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 107 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 107, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1155] = {5'd5, 4'd0, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 107 {'a': 3, 'z': 0, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 107, 'op': 'load'}
    instructions[1156] = {5'd15, 4'd0, 4'd0, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 107 {'a': 0, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 107, 'op': 'write'}
    instructions[1157] = {5'd1, 4'd3, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 107 {'a': 3, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 107, 'op': 'addl'}
    instructions[1158] = {5'd1, 4'd8, 4'd4, 16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108 {'a': 4, 'literal': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108, 'op': 'addl'}
    instructions[1159] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108, 'op': 'addl'}
    instructions[1160] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108, 'op': 'load'}
    instructions[1161] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108, 'op': 'store'}
    instructions[1162] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108, 'op': 'addl'}
    instructions[1163] = {5'd1, 4'd8, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108 {'a': 4, 'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108, 'op': 'addl'}
    instructions[1164] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108, 'op': 'addl'}
    instructions[1165] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108, 'op': 'load'}
    instructions[1166] = {5'd7, 4'd8, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108 {'a': 8, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108, 'op': 'a_lo'}
    instructions[1167] = {5'd8, 4'd0, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108 {'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108, 'op': 'int_to_float'}
    instructions[1168] = {5'd7, 4'd8, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108 {'a': 8, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108, 'op': 'a_lo'}
    instructions[1169] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1170] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108, 'op': 'load'}
    instructions[1171] = {5'd9, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108, 'op': 'float_multiply'}
    instructions[1172] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108, 'op': 'store'}
    instructions[1173] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108, 'op': 'addl'}
    instructions[1174] = {5'd1, 4'd8, 4'd4, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108 {'a': 4, 'literal': -2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108, 'op': 'addl'}
    instructions[1175] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108, 'op': 'addl'}
    instructions[1176] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108, 'op': 'load'}
    instructions[1177] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1178] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108, 'op': 'load'}
    instructions[1179] = {5'd23, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108, 'op': 'float_subtract'}
    instructions[1180] = {5'd1, 4'd2, 4'd4, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108 {'a': 4, 'literal': -2, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108, 'op': 'addl'}
    instructions[1181] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 108, 'op': 'store'}
    instructions[1182] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 109 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 109, 'op': 'literal'}
    instructions[1183] = {5'd6, 4'd8, 4'd8, 16'd16672};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 109 {'a': 8, 'literal': 16672, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 109, 'op': 'literal_hi'}
    instructions[1184] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 109 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 109, 'op': 'store'}
    instructions[1185] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 109 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 109, 'op': 'addl'}
    instructions[1186] = {5'd1, 4'd8, 4'd4, 16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 109 {'a': 4, 'literal': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 109, 'op': 'addl'}
    instructions[1187] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 109 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 109, 'op': 'addl'}
    instructions[1188] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 109 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 109, 'op': 'load'}
    instructions[1189] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 109 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 109, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1190] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 109 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 109, 'op': 'load'}
    instructions[1191] = {5'd24, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 109 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 109, 'op': 'float_divide'}
    instructions[1192] = {5'd1, 4'd2, 4'd4, 16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 109 {'a': 4, 'literal': 2, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 109, 'op': 'addl'}
    instructions[1193] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 109 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 109, 'op': 'store'}
    instructions[1194] = {5'd2, 4'd0, 4'd3, 16'd6};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110, 'op': 'store'}
    instructions[1195] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110, 'op': 'addl'}
    instructions[1196] = {5'd2, 4'd0, 4'd3, 16'd7};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110, 'op': 'store'}
    instructions[1197] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110, 'op': 'addl'}
    instructions[1198] = {5'd1, 4'd8, 4'd4, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110 {'a': 4, 'literal': -2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110, 'op': 'addl'}
    instructions[1199] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110, 'op': 'addl'}
    instructions[1200] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110, 'op': 'load'}
    instructions[1201] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110, 'op': 'store'}
    instructions[1202] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110, 'op': 'addl'}
    instructions[1203] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110, 'op': 'literal'}
    instructions[1204] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110, 'op': 'store'}
    instructions[1205] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110, 'op': 'addl'}
    instructions[1206] = {5'd1, 4'd7, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110 {'a': 4, 'literal': 0, 'z': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110, 'op': 'addl'}
    instructions[1207] = {5'd1, 4'd4, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110 {'a': 3, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110, 'op': 'addl'}
    instructions[1208] = {5'd3, 4'd6, 4'd0, 16'd1414};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110 {'z': 6, 'label': 1414, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110, 'op': 'call'}
    instructions[1209] = {5'd1, 4'd3, 4'd3, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110 {'a': 3, 'literal': -2, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110, 'op': 'addl'}
    instructions[1210] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1211] = {5'd5, 4'd7, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110 {'a': 3, 'z': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110, 'op': 'load'}
    instructions[1212] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1213] = {5'd5, 4'd6, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110 {'a': 3, 'z': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110, 'op': 'load'}
    instructions[1214] = {5'd0, 4'd2, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110 {'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110, 'op': 'literal'}
    instructions[1215] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110, 'op': 'load'}
    instructions[1216] = {5'd14, 4'd0, 4'd8, 16'd1219};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110 {'a': 8, 'label': 1219, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110, 'op': 'jmp_if_false'}
    instructions[1217] = {5'd11, 4'd0, 4'd0, 16'd1222};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110 {'label': 1222, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110, 'op': 'goto'}
    instructions[1218] = {5'd11, 4'd0, 4'd0, 16'd1219};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110 {'label': 1219, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 110, 'op': 'goto'}
    instructions[1219] = {5'd11, 4'd0, 4'd0, 16'd1221};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 112 {'label': 1221, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 112, 'op': 'goto'}
    instructions[1220] = {5'd11, 4'd0, 4'd0, 16'd1222};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 112 {'label': 1222, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 112, 'op': 'goto'}
    instructions[1221] = {5'd11, 4'd0, 4'd0, 16'd1100};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105 {'label': 1100, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 105, 'op': 'goto'}
    instructions[1222] = {5'd1, 4'd3, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 79 {'a': 4, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 79, 'op': 'addl'}
    instructions[1223] = {5'd1, 4'd4, 4'd7, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 79 {'a': 7, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 79, 'op': 'addl'}
    instructions[1224] = {5'd12, 4'd0, 4'd6, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 79 {'a': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/print.h : 79, 'op': 'return'}
    instructions[1225] = {5'd1, 4'd3, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 131 {'a': 3, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 131, 'op': 'addl'}
    instructions[1226] = {5'd1, 4'd8, 4'd4, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 132 {'a': 4, 'literal': -2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 132, 'op': 'addl'}
    instructions[1227] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 132 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 132, 'op': 'addl'}
    instructions[1228] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 132 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 132, 'op': 'load'}
    instructions[1229] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 132 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 132, 'op': 'store'}
    instructions[1230] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 132 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 132, 'op': 'addl'}
    instructions[1231] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 132 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 132, 'op': 'literal'}
    instructions[1232] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 132 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 132, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1233] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 132 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 132, 'op': 'load'}
    instructions[1234] = {5'd26, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 132 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 132, 'op': 'greater'}
    instructions[1235] = {5'd14, 4'd0, 4'd8, 16'd1249};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 132 {'a': 8, 'label': 1249, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 132, 'op': 'jmp_if_false'}
    instructions[1236] = {5'd1, 4'd8, 4'd4, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 133 {'a': 4, 'literal': -2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 133, 'op': 'addl'}
    instructions[1237] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 133 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 133, 'op': 'addl'}
    instructions[1238] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 133 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 133, 'op': 'load'}
    instructions[1239] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 133 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 133, 'op': 'store'}
    instructions[1240] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 133 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 133, 'op': 'addl'}
    instructions[1241] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 133 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 133, 'op': 'literal'}
    instructions[1242] = {5'd6, 4'd8, 4'd8, 16'd32768};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 133 {'a': 8, 'literal': 32768, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 133, 'op': 'literal_hi'}
    instructions[1243] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 133 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 133, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1244] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 133 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 133, 'op': 'load'}
    instructions[1245] = {5'd27, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 133 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 133, 'op': 'subtract'}
    instructions[1246] = {5'd1, 4'd2, 4'd4, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 133 {'a': 4, 'literal': -2, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 133, 'op': 'addl'}
    instructions[1247] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 133 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 133, 'op': 'store'}
    instructions[1248] = {5'd11, 4'd0, 4'd0, 16'd1249};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 132 {'label': 1249, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 132, 'op': 'goto'}
    instructions[1249] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 135 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 135, 'op': 'addl'}
    instructions[1250] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 135 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 135, 'op': 'addl'}
    instructions[1251] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 135 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 135, 'op': 'load'}
    instructions[1252] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 135 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 135, 'op': 'store'}
    instructions[1253] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 135 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 135, 'op': 'addl'}
    instructions[1254] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 135 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 135, 'op': 'literal'}
    instructions[1255] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 135 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 135, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1256] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 135 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 135, 'op': 'load'}
    instructions[1257] = {5'd26, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 135 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 135, 'op': 'greater'}
    instructions[1258] = {5'd14, 4'd0, 4'd8, 16'd1272};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 135 {'a': 8, 'label': 1272, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 135, 'op': 'jmp_if_false'}
    instructions[1259] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 136 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 136, 'op': 'addl'}
    instructions[1260] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 136 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 136, 'op': 'addl'}
    instructions[1261] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 136 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 136, 'op': 'load'}
    instructions[1262] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 136 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 136, 'op': 'store'}
    instructions[1263] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 136 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 136, 'op': 'addl'}
    instructions[1264] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 136 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 136, 'op': 'literal'}
    instructions[1265] = {5'd6, 4'd8, 4'd8, 16'd32768};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 136 {'a': 8, 'literal': 32768, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 136, 'op': 'literal_hi'}
    instructions[1266] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 136 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 136, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1267] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 136 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 136, 'op': 'load'}
    instructions[1268] = {5'd27, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 136 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 136, 'op': 'subtract'}
    instructions[1269] = {5'd1, 4'd2, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 136 {'a': 4, 'literal': -1, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 136, 'op': 'addl'}
    instructions[1270] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 136 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 136, 'op': 'store'}
    instructions[1271] = {5'd11, 4'd0, 4'd0, 16'd1272};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 135 {'label': 1272, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 135, 'op': 'goto'}
    instructions[1272] = {5'd1, 4'd8, 4'd4, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 138 {'a': 4, 'literal': -2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 138, 'op': 'addl'}
    instructions[1273] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 138 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 138, 'op': 'addl'}
    instructions[1274] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 138 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 138, 'op': 'load'}
    instructions[1275] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 138 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 138, 'op': 'store'}
    instructions[1276] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 138 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 138, 'op': 'addl'}
    instructions[1277] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 138 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 138, 'op': 'addl'}
    instructions[1278] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 138 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 138, 'op': 'addl'}
    instructions[1279] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 138 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 138, 'op': 'load'}
    instructions[1280] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 138 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 138, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1281] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 138 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 138, 'op': 'load'}
    instructions[1282] = {5'd26, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 138 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 138, 'op': 'greater'}
    instructions[1283] = {5'd0, 4'd2, 4'd0, 16'd80};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 138 {'literal': 80, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 138, 'op': 'literal'}
    instructions[1284] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 138 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 138, 'op': 'store'}
    instructions[1285] = {5'd1, 4'd3, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 138 {'a': 4, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 138, 'op': 'addl'}
    instructions[1286] = {5'd1, 4'd4, 4'd7, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 138 {'a': 7, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 138, 'op': 'addl'}
    instructions[1287] = {5'd12, 4'd0, 4'd6, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 138 {'a': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 138, 'op': 'return'}
    instructions[1288] = {5'd1, 4'd3, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 161 {'a': 3, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 161, 'op': 'addl'}
    instructions[1289] = {5'd1, 4'd8, 4'd4, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 162 {'a': 4, 'literal': -2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 162, 'op': 'addl'}
    instructions[1290] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 162 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 162, 'op': 'addl'}
    instructions[1291] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 162 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 162, 'op': 'load'}
    instructions[1292] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 162 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 162, 'op': 'store'}
    instructions[1293] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 162 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 162, 'op': 'addl'}
    instructions[1294] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 162 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 162, 'op': 'literal'}
    instructions[1295] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 162 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 162, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1296] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 162 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 162, 'op': 'load'}
    instructions[1297] = {5'd26, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 162 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 162, 'op': 'greater'}
    instructions[1298] = {5'd14, 4'd0, 4'd8, 16'd1312};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 162 {'a': 8, 'label': 1312, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 162, 'op': 'jmp_if_false'}
    instructions[1299] = {5'd1, 4'd8, 4'd4, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 163 {'a': 4, 'literal': -2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 163, 'op': 'addl'}
    instructions[1300] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 163 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 163, 'op': 'addl'}
    instructions[1301] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 163 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 163, 'op': 'load'}
    instructions[1302] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 163 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 163, 'op': 'store'}
    instructions[1303] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 163 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 163, 'op': 'addl'}
    instructions[1304] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 163 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 163, 'op': 'literal'}
    instructions[1305] = {5'd6, 4'd8, 4'd8, 16'd32768};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 163 {'a': 8, 'literal': 32768, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 163, 'op': 'literal_hi'}
    instructions[1306] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 163 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 163, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1307] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 163 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 163, 'op': 'load'}
    instructions[1308] = {5'd27, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 163 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 163, 'op': 'subtract'}
    instructions[1309] = {5'd1, 4'd2, 4'd4, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 163 {'a': 4, 'literal': -2, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 163, 'op': 'addl'}
    instructions[1310] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 163 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 163, 'op': 'store'}
    instructions[1311] = {5'd11, 4'd0, 4'd0, 16'd1312};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 162 {'label': 1312, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 162, 'op': 'goto'}
    instructions[1312] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 165 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 165, 'op': 'addl'}
    instructions[1313] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 165 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 165, 'op': 'addl'}
    instructions[1314] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 165 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 165, 'op': 'load'}
    instructions[1315] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 165 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 165, 'op': 'store'}
    instructions[1316] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 165 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 165, 'op': 'addl'}
    instructions[1317] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 165 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 165, 'op': 'literal'}
    instructions[1318] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 165 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 165, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1319] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 165 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 165, 'op': 'load'}
    instructions[1320] = {5'd26, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 165 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 165, 'op': 'greater'}
    instructions[1321] = {5'd14, 4'd0, 4'd8, 16'd1335};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 165 {'a': 8, 'label': 1335, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 165, 'op': 'jmp_if_false'}
    instructions[1322] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 166 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 166, 'op': 'addl'}
    instructions[1323] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 166 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 166, 'op': 'addl'}
    instructions[1324] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 166 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 166, 'op': 'load'}
    instructions[1325] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 166 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 166, 'op': 'store'}
    instructions[1326] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 166 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 166, 'op': 'addl'}
    instructions[1327] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 166 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 166, 'op': 'literal'}
    instructions[1328] = {5'd6, 4'd8, 4'd8, 16'd32768};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 166 {'a': 8, 'literal': 32768, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 166, 'op': 'literal_hi'}
    instructions[1329] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 166 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 166, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1330] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 166 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 166, 'op': 'load'}
    instructions[1331] = {5'd27, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 166 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 166, 'op': 'subtract'}
    instructions[1332] = {5'd1, 4'd2, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 166 {'a': 4, 'literal': -1, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 166, 'op': 'addl'}
    instructions[1333] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 166 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 166, 'op': 'store'}
    instructions[1334] = {5'd11, 4'd0, 4'd0, 16'd1335};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 165 {'label': 1335, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 165, 'op': 'goto'}
    instructions[1335] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 168 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 168, 'op': 'addl'}
    instructions[1336] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 168 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 168, 'op': 'addl'}
    instructions[1337] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 168 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 168, 'op': 'load'}
    instructions[1338] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 168 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 168, 'op': 'store'}
    instructions[1339] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 168 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 168, 'op': 'addl'}
    instructions[1340] = {5'd1, 4'd8, 4'd4, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 168 {'a': 4, 'literal': -2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 168, 'op': 'addl'}
    instructions[1341] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 168 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 168, 'op': 'addl'}
    instructions[1342] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 168 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 168, 'op': 'load'}
    instructions[1343] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 168 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 168, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1344] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 168 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 168, 'op': 'load'}
    instructions[1345] = {5'd28, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 168 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 168, 'op': 'greater_equal'}
    instructions[1346] = {5'd0, 4'd2, 4'd0, 16'd105};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 168 {'literal': 105, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 168, 'op': 'literal'}
    instructions[1347] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 168 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 168, 'op': 'store'}
    instructions[1348] = {5'd1, 4'd3, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 168 {'a': 4, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 168, 'op': 'addl'}
    instructions[1349] = {5'd1, 4'd4, 4'd7, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 168 {'a': 7, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 168, 'op': 'addl'}
    instructions[1350] = {5'd12, 4'd0, 4'd6, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 168 {'a': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 168, 'op': 'return'}
    instructions[1351] = {5'd1, 4'd3, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 141 {'a': 3, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 141, 'op': 'addl'}
    instructions[1352] = {5'd1, 4'd8, 4'd4, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 142 {'a': 4, 'literal': -2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 142, 'op': 'addl'}
    instructions[1353] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 142 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 142, 'op': 'addl'}
    instructions[1354] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 142 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 142, 'op': 'load'}
    instructions[1355] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 142 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 142, 'op': 'store'}
    instructions[1356] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 142 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 142, 'op': 'addl'}
    instructions[1357] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 142 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 142, 'op': 'literal'}
    instructions[1358] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 142 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 142, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1359] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 142 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 142, 'op': 'load'}
    instructions[1360] = {5'd26, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 142 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 142, 'op': 'greater'}
    instructions[1361] = {5'd14, 4'd0, 4'd8, 16'd1375};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 142 {'a': 8, 'label': 1375, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 142, 'op': 'jmp_if_false'}
    instructions[1362] = {5'd1, 4'd8, 4'd4, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 143 {'a': 4, 'literal': -2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 143, 'op': 'addl'}
    instructions[1363] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 143 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 143, 'op': 'addl'}
    instructions[1364] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 143 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 143, 'op': 'load'}
    instructions[1365] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 143 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 143, 'op': 'store'}
    instructions[1366] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 143 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 143, 'op': 'addl'}
    instructions[1367] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 143 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 143, 'op': 'literal'}
    instructions[1368] = {5'd6, 4'd8, 4'd8, 16'd32768};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 143 {'a': 8, 'literal': 32768, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 143, 'op': 'literal_hi'}
    instructions[1369] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 143 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 143, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1370] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 143 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 143, 'op': 'load'}
    instructions[1371] = {5'd27, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 143 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 143, 'op': 'subtract'}
    instructions[1372] = {5'd1, 4'd2, 4'd4, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 143 {'a': 4, 'literal': -2, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 143, 'op': 'addl'}
    instructions[1373] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 143 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 143, 'op': 'store'}
    instructions[1374] = {5'd11, 4'd0, 4'd0, 16'd1375};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 142 {'label': 1375, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 142, 'op': 'goto'}
    instructions[1375] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 145 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 145, 'op': 'addl'}
    instructions[1376] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 145 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 145, 'op': 'addl'}
    instructions[1377] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 145 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 145, 'op': 'load'}
    instructions[1378] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 145 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 145, 'op': 'store'}
    instructions[1379] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 145 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 145, 'op': 'addl'}
    instructions[1380] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 145 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 145, 'op': 'literal'}
    instructions[1381] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 145 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 145, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1382] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 145 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 145, 'op': 'load'}
    instructions[1383] = {5'd26, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 145 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 145, 'op': 'greater'}
    instructions[1384] = {5'd14, 4'd0, 4'd8, 16'd1398};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 145 {'a': 8, 'label': 1398, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 145, 'op': 'jmp_if_false'}
    instructions[1385] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 146 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 146, 'op': 'addl'}
    instructions[1386] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 146 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 146, 'op': 'addl'}
    instructions[1387] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 146 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 146, 'op': 'load'}
    instructions[1388] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 146 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 146, 'op': 'store'}
    instructions[1389] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 146 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 146, 'op': 'addl'}
    instructions[1390] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 146 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 146, 'op': 'literal'}
    instructions[1391] = {5'd6, 4'd8, 4'd8, 16'd32768};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 146 {'a': 8, 'literal': 32768, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 146, 'op': 'literal_hi'}
    instructions[1392] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 146 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 146, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1393] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 146 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 146, 'op': 'load'}
    instructions[1394] = {5'd27, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 146 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 146, 'op': 'subtract'}
    instructions[1395] = {5'd1, 4'd2, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 146 {'a': 4, 'literal': -1, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 146, 'op': 'addl'}
    instructions[1396] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 146 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 146, 'op': 'store'}
    instructions[1397] = {5'd11, 4'd0, 4'd0, 16'd1398};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 145 {'label': 1398, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 145, 'op': 'goto'}
    instructions[1398] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 148 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 148, 'op': 'addl'}
    instructions[1399] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 148 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 148, 'op': 'addl'}
    instructions[1400] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 148 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 148, 'op': 'load'}
    instructions[1401] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 148 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 148, 'op': 'store'}
    instructions[1402] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 148 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 148, 'op': 'addl'}
    instructions[1403] = {5'd1, 4'd8, 4'd4, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 148 {'a': 4, 'literal': -2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 148, 'op': 'addl'}
    instructions[1404] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 148 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 148, 'op': 'addl'}
    instructions[1405] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 148 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 148, 'op': 'load'}
    instructions[1406] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 148 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 148, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1407] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 148 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 148, 'op': 'load'}
    instructions[1408] = {5'd26, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 148 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 148, 'op': 'greater'}
    instructions[1409] = {5'd0, 4'd2, 4'd0, 16'd82};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 148 {'literal': 82, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 148, 'op': 'literal'}
    instructions[1410] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 148 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 148, 'op': 'store'}
    instructions[1411] = {5'd1, 4'd3, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 148 {'a': 4, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 148, 'op': 'addl'}
    instructions[1412] = {5'd1, 4'd4, 4'd7, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 148 {'a': 7, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 148, 'op': 'addl'}
    instructions[1413] = {5'd12, 4'd0, 4'd6, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 148 {'a': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 148, 'op': 'return'}
    instructions[1414] = {5'd1, 4'd3, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 111 {'a': 3, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 111, 'op': 'addl'}
    instructions[1415] = {5'd1, 4'd8, 4'd4, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 112 {'a': 4, 'literal': -2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 112, 'op': 'addl'}
    instructions[1416] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 112 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 112, 'op': 'addl'}
    instructions[1417] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 112 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 112, 'op': 'load'}
    instructions[1418] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 112 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 112, 'op': 'store'}
    instructions[1419] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 112 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 112, 'op': 'addl'}
    instructions[1420] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 112 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 112, 'op': 'literal'}
    instructions[1421] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 112 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 112, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1422] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 112 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 112, 'op': 'load'}
    instructions[1423] = {5'd26, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 112 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 112, 'op': 'greater'}
    instructions[1424] = {5'd14, 4'd0, 4'd8, 16'd1438};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 112 {'a': 8, 'label': 1438, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 112, 'op': 'jmp_if_false'}
    instructions[1425] = {5'd1, 4'd8, 4'd4, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 113 {'a': 4, 'literal': -2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 113, 'op': 'addl'}
    instructions[1426] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 113 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 113, 'op': 'addl'}
    instructions[1427] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 113 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 113, 'op': 'load'}
    instructions[1428] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 113 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 113, 'op': 'store'}
    instructions[1429] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 113 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 113, 'op': 'addl'}
    instructions[1430] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 113 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 113, 'op': 'literal'}
    instructions[1431] = {5'd6, 4'd8, 4'd8, 16'd32768};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 113 {'a': 8, 'literal': 32768, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 113, 'op': 'literal_hi'}
    instructions[1432] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 113 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 113, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1433] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 113 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 113, 'op': 'load'}
    instructions[1434] = {5'd27, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 113 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 113, 'op': 'subtract'}
    instructions[1435] = {5'd1, 4'd2, 4'd4, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 113 {'a': 4, 'literal': -2, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 113, 'op': 'addl'}
    instructions[1436] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 113 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 113, 'op': 'store'}
    instructions[1437] = {5'd11, 4'd0, 4'd0, 16'd1438};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 112 {'label': 1438, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 112, 'op': 'goto'}
    instructions[1438] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 115 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 115, 'op': 'addl'}
    instructions[1439] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 115 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 115, 'op': 'addl'}
    instructions[1440] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 115 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 115, 'op': 'load'}
    instructions[1441] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 115 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 115, 'op': 'store'}
    instructions[1442] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 115 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 115, 'op': 'addl'}
    instructions[1443] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 115 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 115, 'op': 'literal'}
    instructions[1444] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 115 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 115, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1445] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 115 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 115, 'op': 'load'}
    instructions[1446] = {5'd26, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 115 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 115, 'op': 'greater'}
    instructions[1447] = {5'd14, 4'd0, 4'd8, 16'd1461};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 115 {'a': 8, 'label': 1461, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 115, 'op': 'jmp_if_false'}
    instructions[1448] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 116 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 116, 'op': 'addl'}
    instructions[1449] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 116 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 116, 'op': 'addl'}
    instructions[1450] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 116 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 116, 'op': 'load'}
    instructions[1451] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 116 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 116, 'op': 'store'}
    instructions[1452] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 116 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 116, 'op': 'addl'}
    instructions[1453] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 116 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 116, 'op': 'literal'}
    instructions[1454] = {5'd6, 4'd8, 4'd8, 16'd32768};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 116 {'a': 8, 'literal': 32768, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 116, 'op': 'literal_hi'}
    instructions[1455] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 116 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 116, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1456] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 116 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 116, 'op': 'load'}
    instructions[1457] = {5'd27, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 116 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 116, 'op': 'subtract'}
    instructions[1458] = {5'd1, 4'd2, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 116 {'a': 4, 'literal': -1, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 116, 'op': 'addl'}
    instructions[1459] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 116 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 116, 'op': 'store'}
    instructions[1460] = {5'd11, 4'd0, 4'd0, 16'd1461};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 115 {'label': 1461, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 115, 'op': 'goto'}
    instructions[1461] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 118 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 118, 'op': 'addl'}
    instructions[1462] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 118 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 118, 'op': 'addl'}
    instructions[1463] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 118 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 118, 'op': 'load'}
    instructions[1464] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 118 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 118, 'op': 'store'}
    instructions[1465] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 118 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 118, 'op': 'addl'}
    instructions[1466] = {5'd1, 4'd8, 4'd4, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 118 {'a': 4, 'literal': -2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 118, 'op': 'addl'}
    instructions[1467] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 118 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 118, 'op': 'addl'}
    instructions[1468] = {5'd5, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 118 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 118, 'op': 'load'}
    instructions[1469] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 118 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 118, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[1470] = {5'd5, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 118 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 118, 'op': 'load'}
    instructions[1471] = {5'd29, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 118 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 118, 'op': 'equal'}
    instructions[1472] = {5'd0, 4'd2, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 118 {'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 118, 'op': 'literal'}
    instructions[1473] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 118 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 118, 'op': 'store'}
    instructions[1474] = {5'd1, 4'd3, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 118 {'a': 4, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 118, 'op': 'addl'}
    instructions[1475] = {5'd1, 4'd4, 4'd7, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 118 {'a': 7, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 118, 'op': 'addl'}
    instructions[1476] = {5'd12, 4'd0, 4'd6, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 118 {'a': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/builtins.h : 118, 'op': 'return'}
  end

  
  always @(posedge clk)
  begin
    load_data <= memory[load_address];
    if(store_enable && state == execute) begin
      memory[store_address] <= store_data;
    end
  end


  //////////////////////////////////////////////////////////////////////////////
  // PIPELINE STAGE 1 -- FETCH INSTRUCTION
  //                                                                            
  
  always @(posedge clk)
  begin
    //implement memory for instructions
    if (state == instruction_fetch || state == operand_fetch || state == execute) begin
      instruction <= instructions[program_counter];
      program_counter_1 <= program_counter;
    end
  end

  assign opcode    = instruction[28:24];
  assign address_z = instruction[23:20];
  assign address_a = instruction[19:16];
  assign address_b = instruction[3:0];
  assign literal   = instruction[15:0];

  //////////////////////////////////////////////////////////////////////////////
  // PIPELINE STAGE 2 -- FETCH OPERANDS
  //                                                                            
  
  always @(posedge clk)
  begin
    if (write_enable) begin
      registers[address_z_3] <= result;
    end
    if (state == operand_fetch || state == execute) begin
      opcode_2 <= opcode;
      literal_2 <= literal;
      address_a_2 <= address_a;
      address_b_2 <= address_b;
      address_z_2 <= address_z;
      program_counter_2 <= program_counter_1;
    end
  end
  assign register_a = registers[address_a_2];
  assign register_b = registers[address_b_2];
  assign operand_a = (address_a_2 == address_z_3 && write_enable)?result:register_a;
  assign operand_b = (address_b_2 == address_z_3 && write_enable)?result:register_b;
  assign store_address = operand_a;
  assign load_address = operand_a;
  assign store_data = operand_b;
  assign store_enable = (opcode_2==2);

  //////////////////////////////////////////////////////////////////////////////
  // PIPELINE STAGE 3 -- EXECUTE
  //                                                                            
  
  always @(posedge clk)
  begin

  write_enable <= 0;
  timer_clock <= timer_clock + 1;
  case(state)

    //instruction_fetch
    instruction_fetch: begin
      program_counter <= program_counter + 1;
      state <= operand_fetch;
    end
    //operand_fetch
    operand_fetch: begin
      program_counter <= program_counter + 1;
      state <= execute;
    end
    //execute
    execute: begin
      program_counter <= program_counter + 1;
      address_z_3 <= address_z_2;
      case(opcode_2)

        //literal
        16'd0:
        begin
          result<=$signed(literal_2);
          write_enable <= 1;
        end

        //addl
        16'd1:
        begin
          result<=operand_a + literal_2;
          write_enable <= 1;
        end

        //store
        16'd2:
        begin
        end

        //call
        16'd3:
        begin
          result <= program_counter_2 + 1;
          write_enable <= 1;
          program_counter <= literal_2;
          state <= instruction_fetch;
        end

        //stop
        16'd4:
        begin
        state <= stop;
        end

        //load
        16'd5:
        begin
          state <= load;
        end

        //literal_hi
        16'd6:
        begin
          result<= {literal_2, operand_a[15:0]};
          write_enable <= 1;
        end

        //a_lo
        16'd7:
        begin
          a_lo <= operand_a;
          result <= a_lo;
          write_enable <= 1;
        end

        //int_to_float
        16'd8:
        begin
          int_to_float_in <= a_lo;
          state <= int_to_float_write_a;
        end

        //float_multiply
        16'd9:
        begin
          multiplier_a_stb <= 1;
          multiplier_a <= operand_a;
          multiplier_b <= operand_b;
          state <= multiplier_write_a;
        end

        //wait_clocks
        16'd10:
        begin
          timer <= operand_a;
          state <= wait_state;
        end

        //goto
        16'd11:
        begin
          program_counter <= literal_2;
          state <= instruction_fetch;
        end

        //return
        16'd12:
        begin
          program_counter <= operand_a;
          state <= instruction_fetch;
        end

        //add
        16'd13:
        begin
          long_result = operand_a + operand_b;
          result <= long_result[31:0];
          carry[0] <= long_result[32];
          write_enable <= 1;
        end

        //jmp_if_false
        16'd14:
        begin
          if (operand_a == 0) begin
            program_counter <= literal_2;
            state <= instruction_fetch;
          end
        end

        //write
        16'd15:
        begin
          state <= write;
          write_output <= operand_a;
          write_value <= operand_b;
        end

        //timer_low
        16'd16:
        begin
          result <= timer_clock[31:0];
          write_enable <= 1;
        end

        //unsigned_greater
        16'd17:
        begin
          result <= $unsigned(operand_a) > $unsigned(operand_b);
          write_enable <= 1;
        end

        //or
        16'd18:
        begin
          result <= operand_a | operand_b;
          write_enable <= 1;
        end

        //shift_left
        16'd19:
        begin
          if(operand_b < 32) begin
            result <= operand_a << operand_b;
            carry <= operand_a >> (32-operand_b);
          end else begin
            result <= 0;
            carry <= operand_a;
          end
          write_enable <= 1;
        end

        //unsigned_shift_right
        16'd20:
        begin
          if(operand_b < 32) begin
            result <= operand_a >> operand_b;
            carry <= operand_a << (32-operand_b);
          end else begin
            result <= 0;
            carry <= operand_a;
          end
          write_enable <= 1;
        end

        //read
        16'd21:
        begin
          state <= read;
          read_input <= operand_a;
        end

        //and
        16'd22:
        begin
          result <= operand_a & operand_b;
          write_enable <= 1;
        end

        //float_subtract
        16'd23:
        begin
          adder_a_stb <= 1;
          adder_a <= operand_a;
          adder_b <= {~operand_b[31], operand_b[30:0]};
          state <= adder_write_a;
        end

        //float_divide
        16'd24:
        begin
          divider_a_stb <= 1;
          divider_a <= operand_a;
          divider_b <= operand_b;
          state <= divider_write_a;
        end

        //float_to_int
        16'd25:
        begin
          float_to_int_in <= a_lo;
          state <= float_to_int_write_a;
        end

        //greater
        16'd26:
        begin
          result <= $signed(operand_a) > $signed(operand_b);
          write_enable <= 1;
        end

        //subtract
        16'd27:
        begin
          long_result = operand_a + (~operand_b) + 1;
          result <= long_result[31:0];
          carry[0] <= ~long_result[32];
          write_enable <= 1;
        end

        //greater_equal
        16'd28:
        begin
          result <= $signed(operand_a) >= $signed(operand_b);
          write_enable <= 1;
        end

        //equal
        16'd29:
        begin
          result <= operand_a == operand_b;
          write_enable <= 1;
        end

      endcase

    end

    read:
    begin
      case(read_input)
      0:
      begin
        s_input_i2c_in_ack <= 1;
        if (s_input_i2c_in_ack && input_i2c_in_stb) begin
          result <= input_i2c_in;
          write_enable <= 1;
          s_input_i2c_in_ack <= 0;
          state <= execute;
        end
      end
      endcase
    end

    write:
    begin
      case(write_output)
      1:
      begin
        s_output_i2c_out_stb <= 1;
        s_output_i2c_out <= write_value;
        if (output_i2c_out_ack && s_output_i2c_out_stb) begin
          s_output_i2c_out_stb <= 0;
          state <= execute;
        end
      end
      2:
      begin
        s_output_rs232_tx_stb <= 1;
        s_output_rs232_tx <= write_value;
        if (output_rs232_tx_ack && s_output_rs232_tx_stb) begin
          s_output_rs232_tx_stb <= 0;
          state <= execute;
        end
      end
      endcase
    end

    load:
    begin
        result <= load_data;
        write_enable <= 1;
        state <= execute;
    end

    wait_state:
    begin
      if (timer) begin
        timer <= timer - 1;
      end else begin
        state <= execute;
      end
    end

    stop:
    begin
    end

    divider_write_a:
    begin
      divider_a_stb <= 1;
      if (divider_a_stb && divider_a_ack) begin
        divider_a_stb <= 0;
        state <= divider_write_b;
      end
    end

    divider_write_b:
    begin
      divider_b_stb <= 1;
      if (divider_b_stb && divider_b_ack) begin
        divider_b_stb <= 0;
        state <= divider_read_z;
      end
    end

    divider_read_z:
    begin
      divider_z_ack <= 1;
      if (divider_z_stb && divider_z_ack) begin
        result <= divider_z;
        write_enable <= 1;
        divider_z_ack <= 0;
        state <= execute;
      end
    end

    adder_write_a:
    begin
      adder_a_stb <= 1;
      if (adder_a_stb && adder_a_ack) begin
        adder_a_stb <= 0;
        state <= adder_write_b;
      end
    end

    adder_write_b:
    begin
      adder_b_stb <= 1;
      if (adder_b_stb && adder_b_ack) begin
        adder_b_stb <= 0;
        state <= adder_read_z;
      end
    end

    adder_read_z:
    begin
      adder_z_ack <= 1;
      if (adder_z_stb && adder_z_ack) begin
        result <= adder_z;
        write_enable <= 1;
        adder_z_ack <= 0;
        state <= execute;
      end
    end

    multiplier_write_a:
    begin
      multiplier_a_stb <= 1;
      if (multiplier_a_stb && multiplier_a_ack) begin
        multiplier_a_stb <= 0;
        state <= multiplier_write_b;
      end
    end

    multiplier_write_b:
    begin
      multiplier_b_stb <= 1;
      if (multiplier_b_stb && multiplier_b_ack) begin
        multiplier_b_stb <= 0;
        state <= multiplier_read_z;
      end
    end

    multiplier_read_z:
    begin
      multiplier_z_ack <= 1;
      if (multiplier_z_stb && multiplier_z_ack) begin
        result <= multiplier_z;
        write_enable <= 1;
        multiplier_z_ack <= 0;
        state <= execute;
      end
    end

     int_to_float_write_a:
     begin
       int_to_float_in_stb <= 1;
       if (int_to_float_in_stb && int_to_float_in_ack) begin
         int_to_float_in_stb <= 0;
         state <= int_to_float_read_z;
       end
     end

     int_to_float_read_z:
     begin
       int_to_float_out_ack <= 1;
       if (int_to_float_out_stb && int_to_float_out_ack) begin
         int_to_float_out_ack <= 0;
         a_lo <= int_to_float_out;
         state <= execute;
       end
     end

     float_to_int_write_a:
     begin
       float_to_int_in_stb <= 1;
       if (float_to_int_in_stb && float_to_int_in_ack) begin
         float_to_int_in_stb <= 0;
         state <= float_to_int_read_z;
       end
     end

     float_to_int_read_z:
     begin
       float_to_int_out_ack <= 1;
       if (float_to_int_out_stb && float_to_int_out_ack) begin
         float_to_int_out_ack <= 0;
         a_lo <= float_to_int_out;
         state <= execute;
       end
     end

    endcase

    if (rst == 1'b1) begin
      timer <= 0;
      timer_clock <= 0;
      program_counter <= 0;
      address_z_3 <= 0;
      result <= 0;
      a = 0;
      b = 0;
      z = 0;
      state <= instruction_fetch;
      s_input_i2c_in_ack <= 0;
      s_output_i2c_out_stb <= 0;
      s_output_rs232_tx_stb <= 0;
      divider_a_stb <= 0;
      divider_b_stb <= 0;
      divider_z_ack <= 0;
      adder_a_stb <= 0;
      adder_b_stb <= 0;
      adder_z_ack <= 0;
      multiplier_a_stb <= 0;
      multiplier_b_stb <= 0;
      multiplier_z_ack <= 0;
      int_to_float_in_stb <= 0;
      int_to_float_out_ack <= 0;
      float_to_int_in_stb <= 0;
      float_to_int_out_ack <= 0;
    end
  end
  assign input_i2c_in_ack = s_input_i2c_in_ack;
  assign output_i2c_out_stb = s_output_i2c_out_stb;
  assign output_i2c_out = s_output_i2c_out;
  assign output_rs232_tx_stb = s_output_rs232_tx_stb;
  assign output_rs232_tx = s_output_rs232_tx;

endmodule
