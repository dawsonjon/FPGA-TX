//name : main_0
//input : input_eth_in:16
//input : input_audio_in:16
//input : input_rs232_rx:16
//output : output_eth_out:16
//output : output_audio_out:16
//output : output_frequency_out:16
//output : output_samples_out:16
//output : output_rs232_tx:16
//source_file : /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c

///+============================================================================+
///|                                                                            |
///|                     This file was generated by Chips                       |
///|                                                                            |
///|                                  Chips                                     |
///|                                                                            |
///|                      http://github.com/dawsonjon/Chips-2.0                 |
///|                                                                            |
///|                                                             Python powered |
///+============================================================================+
module main_0(input_eth_in,input_audio_in,input_rs232_rx,input_eth_in_stb,input_audio_in_stb,input_rs232_rx_stb,output_eth_out_ack,output_audio_out_ack,output_frequency_out_ack,output_samples_out_ack,output_rs232_tx_ack,clk,rst,output_eth_out,output_audio_out,output_frequency_out,output_samples_out,output_rs232_tx,output_eth_out_stb,output_audio_out_stb,output_frequency_out_stb,output_samples_out_stb,output_rs232_tx_stb,input_eth_in_ack,input_audio_in_ack,input_rs232_rx_ack,exception);
  integer file_count;
  reg [63:0] double_divider_a;
  reg [63:0] double_divider_b;
  wire [63:0] double_divider_z;
  reg double_divider_a_stb;
  wire double_divider_a_ack;
  reg double_divider_b_stb;
  wire double_divider_b_ack;
  wire double_divider_z_stb;
  reg double_divider_z_ack;
  reg [63:0] double_to_long_in;
  wire [63:0] double_to_long_out;
  wire double_to_long_out_stb;
  reg double_to_long_out_ack;
  reg double_to_long_in_stb;
  wire double_to_long_in_ack;
  reg [63:0] long_to_double_in;
  wire [63:0] long_to_double_out;
  wire long_to_double_out_stb;
  reg long_to_double_out_ack;
  reg long_to_double_in_stb;
  wire long_to_double_in_ack;
  parameter  stop = 4'd0,
  instruction_fetch = 4'd1,
  operand_fetch = 4'd2,
  execute = 4'd3,
  load = 4'd4,
  wait_state = 4'd5,
  read = 4'd6,
  write = 4'd7,
  multiply = 4'd8,
  double_divider_write_a = 4'd9,
  double_divider_write_b = 4'd10,
  double_divider_read_z = 4'd11,
  double_to_long_write_a = 4'd12,
  double_to_long_read_z = 4'd13,
  long_to_double_write_a = 4'd14,
  long_to_double_read_z = 4'd15;
  input [31:0] input_eth_in;
  input [31:0] input_audio_in;
  input [31:0] input_rs232_rx;
  input input_eth_in_stb;
  input input_audio_in_stb;
  input input_rs232_rx_stb;
  input output_eth_out_ack;
  input output_audio_out_ack;
  input output_frequency_out_ack;
  input output_samples_out_ack;
  input output_rs232_tx_ack;
  input clk;
  input rst;
  output [31:0] output_eth_out;
  output [31:0] output_audio_out;
  output [31:0] output_frequency_out;
  output [31:0] output_samples_out;
  output [31:0] output_rs232_tx;
  output output_eth_out_stb;
  output output_audio_out_stb;
  output output_frequency_out_stb;
  output output_samples_out_stb;
  output output_rs232_tx_stb;
  output input_eth_in_ack;
  output input_audio_in_ack;
  output input_rs232_rx_ack;
  reg [31:0] timer;
  reg [63:0] timer_clock;
  reg [15:0] program_counter;
  reg [15:0] program_counter_1;
  reg [15:0] program_counter_2;
  reg [44:0] instruction;
  reg [4:0] opcode_2;
  reg [3:0] a;
  reg [3:0] b;
  reg [3:0] z;
  reg write_enable;
  reg [3:0] address_a_2;
  reg [3:0] address_b_2;
  reg [3:0] address_z_2;
  reg [3:0] address_z_3;
  reg [31:0] load_data;
  reg [31:0] write_output;
  reg [31:0] write_value;
  reg [31:0] read_input;
  reg [15:0] literal_2;
  reg [31:0] a_hi;
  reg [31:0] b_hi;
  reg [31:0] a_lo;
  reg [31:0] b_lo;
  reg [63:0] long_result;
  reg [31:0] result;
  reg [15:0] address;
  reg [31:0] data_out;
  reg [31:0] data_in;
  reg [31:0] carry;
  reg [31:0] s_output_eth_out_stb;
  reg [31:0] s_output_audio_out_stb;
  reg [31:0] s_output_frequency_out_stb;
  reg [31:0] s_output_samples_out_stb;
  reg [31:0] s_output_rs232_tx_stb;
  reg [31:0] s_output_eth_out;
  reg [31:0] s_output_audio_out;
  reg [31:0] s_output_frequency_out;
  reg [31:0] s_output_samples_out;
  reg [31:0] s_output_rs232_tx;
  reg [31:0] s_input_eth_in_ack;
  reg [31:0] s_input_audio_in_ack;
  reg [31:0] s_input_rs232_rx_ack;
  reg [15:0] state;
  output reg exception;
  reg [28:0] instructions [922:0];
  reg [31:0] memory [4096:0];
  reg [31:0] registers [15:0];
  wire [31:0] operand_a;
  wire [31:0] operand_b;
  wire [31:0] register_a;
  wire [31:0] register_b;
  wire [15:0] literal;
  wire [4:0] opcode;
  wire [3:0] address_a;
  wire [3:0] address_b;
  wire [3:0] address_z;
  wire [15:0] load_address;
  wire [15:0] store_address;
  wire [31:0] store_data;
  wire  store_enable;
  reg [31:0] product_a;
  reg [31:0] product_b;
  reg [31:0] product_c;
  reg [31:0] product_d;

  //////////////////////////////////////////////////////////////////////////////
  // Floating Point Arithmetic                                                  
  //                                                                            
  // Generate IEEE 754 single precision divider, adder and multiplier           
  //                                                                            
  double_divider double_divider_inst(
    .clk(clk),
    .rst(rst),
    .input_a(double_divider_a),
    .input_a_stb(double_divider_a_stb),
    .input_a_ack(double_divider_a_ack),
    .input_b(double_divider_b),
    .input_b_stb(double_divider_b_stb),
    .input_b_ack(double_divider_b_ack),
    .output_z(double_divider_z),
    .output_z_stb(double_divider_z_stb),
    .output_z_ack(double_divider_z_ack)
  );
  double_to_long double_to_long_inst(
    .clk(clk),
    .rst(rst),
    .input_a(double_to_long_in),
    .input_a_stb(double_to_long_in_stb),
    .input_a_ack(double_to_long_in_ack),
    .output_z(double_to_long_out),
    .output_z_stb(double_to_long_out_stb),
    .output_z_ack(double_to_long_out_ack)
  );
  long_to_double long_to_double_inst(
    .clk(clk),
    .rst(rst),
    .input_a(long_to_double_in),
    .input_a_stb(long_to_double_in_stb),
    .input_a_ack(long_to_double_in_ack),
    .output_z(long_to_double_out),
    .output_z_stb(long_to_double_out_stb),
    .output_z_ack(long_to_double_out_ack)
  );

  //////////////////////////////////////////////////////////////////////////////
  // INSTRUCTION INITIALIZATION                                                 
  //                                                                            
  // Initialise the contents of the instruction memory                          
  //
  // Intruction Set
  // ==============
  // 0 {'literal': True, 'op': 'literal'}
  // 1 {'literal': True, 'op': 'addl'}
  // 2 {'literal': False, 'op': 'store'}
  // 3 {'literal': True, 'op': 'call'}
  // 4 {'literal': False, 'op': 'stop'}
  // 5 {'literal': True, 'op': 'literal_hi'}
  // 6 {'literal': False, 'op': 'load'}
  // 7 {'literal': False, 'op': 'write'}
  // 8 {'literal': False, 'op': 'a_hi'}
  // 9 {'literal': False, 'op': 'a_lo'}
  // 10 {'literal': False, 'op': 'long_to_double'}
  // 11 {'literal': False, 'op': 'b_hi'}
  // 12 {'literal': False, 'op': 'b_lo'}
  // 13 {'literal': False, 'op': 'long_float_divide'}
  // 14 {'literal': False, 'op': 'double_to_long'}
  // 15 {'literal': False, 'op': 'read'}
  // 16 {'literal': False, 'op': 'shift_right'}
  // 17 {'literal': False, 'op': 'subtract'}
  // 18 {'literal': False, 'op': 'add'}
  // 19 {'literal': False, 'op': 'greater'}
  // 20 {'literal': True, 'op': 'jmp_if_false'}
  // 21 {'literal': True, 'op': 'goto'}
  // 22 {'literal': False, 'op': 'equal'}
  // 23 {'literal': False, 'op': 'return'}
  // 24 {'literal': False, 'op': 'multiply'}
  // 25 {'literal': False, 'op': 'greater_equal'}
  // Intructions
  // ===========
  
  initial
  begin
    instructions[0] = {5'd0, 4'd3, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 94 {'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 94, 'op': 'literal'}
    instructions[1] = {5'd0, 4'd4, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 94 {'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 94, 'op': 'literal'}
    instructions[2] = {5'd1, 4'd3, 4'd3, 16'd75};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 94 {'a': 3, 'literal': 75, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 94, 'op': 'addl'}
    instructions[3] = {5'd0, 4'd8, 4'd0, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 7 {'literal': 4, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 7, 'op': 'literal'}
    instructions[4] = {5'd0, 4'd2, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 7 {'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 7, 'op': 'literal'}
    instructions[5] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 7 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 7, 'op': 'store'}
    instructions[6] = {5'd0, 4'd8, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 4 {'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 4, 'op': 'literal'}
    instructions[7] = {5'd0, 4'd2, 4'd0, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 4 {'literal': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 4, 'op': 'literal'}
    instructions[8] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 4 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 4, 'op': 'store'}
    instructions[9] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 5 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 5, 'op': 'literal'}
    instructions[10] = {5'd0, 4'd2, 4'd0, 16'd4};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 5 {'literal': 4, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 5, 'op': 'literal'}
    instructions[11] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 5 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 5, 'op': 'store'}
    instructions[12] = {5'd0, 4'd8, 4'd0, 16'd5};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 8 {'literal': 5, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 8, 'op': 'literal'}
    instructions[13] = {5'd0, 4'd2, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 8 {'literal': 6, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 8, 'op': 'literal'}
    instructions[14] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 8 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 8, 'op': 'store'}
    instructions[15] = {5'd0, 4'd8, 4'd0, 16'd99};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 99, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[16] = {5'd0, 4'd2, 4'd0, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 7, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[17] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'store'}
    instructions[18] = {5'd0, 4'd8, 4'd0, 16'd97};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 97, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[19] = {5'd0, 4'd2, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 8, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[20] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'store'}
    instructions[21] = {5'd0, 4'd8, 4'd0, 16'd108};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 108, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[22] = {5'd0, 4'd2, 4'd0, 16'd9};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 9, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[23] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'store'}
    instructions[24] = {5'd0, 4'd8, 4'd0, 16'd99};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 99, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[25] = {5'd0, 4'd2, 4'd0, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 10, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[26] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'store'}
    instructions[27] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[28] = {5'd0, 4'd2, 4'd0, 16'd11};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 11, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[29] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'store'}
    instructions[30] = {5'd0, 4'd8, 4'd0, 16'd108};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 108, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[31] = {5'd0, 4'd2, 4'd0, 16'd12};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 12, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[32] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'store'}
    instructions[33] = {5'd0, 4'd8, 4'd0, 16'd97};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 97, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[34] = {5'd0, 4'd2, 4'd0, 16'd13};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 13, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[35] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'store'}
    instructions[36] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[37] = {5'd0, 4'd2, 4'd0, 16'd14};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 14, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[38] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'store'}
    instructions[39] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[40] = {5'd0, 4'd2, 4'd0, 16'd15};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 15, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[41] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'store'}
    instructions[42] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[43] = {5'd0, 4'd2, 4'd0, 16'd16};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 16, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[44] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'store'}
    instructions[45] = {5'd0, 4'd8, 4'd0, 16'd103};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 103, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[46] = {5'd0, 4'd2, 4'd0, 16'd17};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 17, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[47] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'store'}
    instructions[48] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[49] = {5'd0, 4'd2, 4'd0, 16'd18};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 18, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[50] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'store'}
    instructions[51] = {5'd0, 4'd8, 4'd0, 16'd102};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 102, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[52] = {5'd0, 4'd2, 4'd0, 16'd19};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 19, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[53] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'store'}
    instructions[54] = {5'd0, 4'd8, 4'd0, 16'd114};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 114, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[55] = {5'd0, 4'd2, 4'd0, 16'd20};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 20, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[56] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'store'}
    instructions[57] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[58] = {5'd0, 4'd2, 4'd0, 16'd21};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 21, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[59] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'store'}
    instructions[60] = {5'd0, 4'd8, 4'd0, 16'd113};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 113, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[61] = {5'd0, 4'd2, 4'd0, 16'd22};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 22, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[62] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'store'}
    instructions[63] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[64] = {5'd0, 4'd2, 4'd0, 16'd23};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 23, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[65] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'store'}
    instructions[66] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[67] = {5'd0, 4'd2, 4'd0, 16'd24};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 24, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[68] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'store'}
    instructions[69] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[70] = {5'd0, 4'd2, 4'd0, 16'd25};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 25, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[71] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'store'}
    instructions[72] = {5'd0, 4'd8, 4'd0, 16'd99};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 99, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[73] = {5'd0, 4'd2, 4'd0, 16'd26};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 26, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[74] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'store'}
    instructions[75] = {5'd0, 4'd8, 4'd0, 16'd121};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 121, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[76] = {5'd0, 4'd2, 4'd0, 16'd27};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 27, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[77] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'store'}
    instructions[78] = {5'd0, 4'd8, 4'd0, 16'd58};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 58, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[79] = {5'd0, 4'd2, 4'd0, 16'd28};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 28, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[80] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'store'}
    instructions[81] = {5'd0, 4'd8, 4'd0, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 10, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[82] = {5'd0, 4'd2, 4'd0, 16'd29};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 29, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[83] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'store'}
    instructions[84] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[85] = {5'd0, 4'd2, 4'd0, 16'd30};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 30, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[86] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'store'}
    instructions[87] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 4 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 4, 'op': 'literal'}
    instructions[88] = {5'd0, 4'd2, 4'd0, 16'd31};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 4 {'literal': 31, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 4, 'op': 'literal'}
    instructions[89] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 4 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 4, 'op': 'store'}
    instructions[90] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 3 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 3, 'op': 'literal'}
    instructions[91] = {5'd0, 4'd2, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 3 {'literal': 32, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 3, 'op': 'literal'}
    instructions[92] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 3 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 3, 'op': 'store'}
    instructions[93] = {5'd0, 4'd8, 4'd0, 16'd69};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 69, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[94] = {5'd0, 4'd2, 4'd0, 16'd33};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 33, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[95] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'store'}
    instructions[96] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[97] = {5'd0, 4'd2, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 34, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[98] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'store'}
    instructions[99] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[100] = {5'd0, 4'd2, 4'd0, 16'd35};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 35, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[101] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'store'}
    instructions[102] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[103] = {5'd0, 4'd2, 4'd0, 16'd36};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 36, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[104] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'store'}
    instructions[105] = {5'd0, 4'd8, 4'd0, 16'd114};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 114, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[106] = {5'd0, 4'd2, 4'd0, 16'd37};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 37, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[107] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'store'}
    instructions[108] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[109] = {5'd0, 4'd2, 4'd0, 16'd38};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 38, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[110] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'store'}
    instructions[111] = {5'd0, 4'd8, 4'd0, 16'd102};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 102, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[112] = {5'd0, 4'd2, 4'd0, 16'd39};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 39, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[113] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'store'}
    instructions[114] = {5'd0, 4'd8, 4'd0, 16'd114};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 114, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[115] = {5'd0, 4'd2, 4'd0, 16'd40};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 40, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[116] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'store'}
    instructions[117] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[118] = {5'd0, 4'd2, 4'd0, 16'd41};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 41, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[119] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'store'}
    instructions[120] = {5'd0, 4'd8, 4'd0, 16'd113};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 113, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[121] = {5'd0, 4'd2, 4'd0, 16'd42};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 42, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[122] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'store'}
    instructions[123] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[124] = {5'd0, 4'd2, 4'd0, 16'd43};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 43, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[125] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'store'}
    instructions[126] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[127] = {5'd0, 4'd2, 4'd0, 16'd44};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 44, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[128] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'store'}
    instructions[129] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[130] = {5'd0, 4'd2, 4'd0, 16'd45};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 45, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[131] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'store'}
    instructions[132] = {5'd0, 4'd8, 4'd0, 16'd99};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 99, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[133] = {5'd0, 4'd2, 4'd0, 16'd46};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 46, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[134] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'store'}
    instructions[135] = {5'd0, 4'd8, 4'd0, 16'd121};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 121, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[136] = {5'd0, 4'd2, 4'd0, 16'd47};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 47, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[137] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'store'}
    instructions[138] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[139] = {5'd0, 4'd2, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 48, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[140] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'store'}
    instructions[141] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[142] = {5'd0, 4'd2, 4'd0, 16'd49};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 49, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[143] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'store'}
    instructions[144] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[145] = {5'd0, 4'd2, 4'd0, 16'd50};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 50, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[146] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'store'}
    instructions[147] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[148] = {5'd0, 4'd2, 4'd0, 16'd51};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 51, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[149] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'store'}
    instructions[150] = {5'd0, 4'd8, 4'd0, 16'd104};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 104, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[151] = {5'd0, 4'd2, 4'd0, 16'd52};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 52, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[152] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'store'}
    instructions[153] = {5'd0, 4'd8, 4'd0, 16'd122};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 122, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[154] = {5'd0, 4'd2, 4'd0, 16'd53};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 53, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[155] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'store'}
    instructions[156] = {5'd0, 4'd8, 4'd0, 16'd58};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 58, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[157] = {5'd0, 4'd2, 4'd0, 16'd54};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 54, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[158] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'store'}
    instructions[159] = {5'd0, 4'd8, 4'd0, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 10, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[160] = {5'd0, 4'd2, 4'd0, 16'd55};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 55, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[161] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'store'}
    instructions[162] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[163] = {5'd0, 4'd2, 4'd0, 16'd56};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 56, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[164] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'store'}
    instructions[165] = {5'd0, 4'd8, 4'd0, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 10 {'literal': 7, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 10, 'op': 'literal'}
    instructions[166] = {5'd0, 4'd2, 4'd0, 16'd57};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 10 {'literal': 57, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 10, 'op': 'literal'}
    instructions[167] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 10 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 10, 'op': 'store'}
    instructions[168] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'literal'}
    instructions[169] = {5'd0, 4'd2, 4'd0, 16'd58};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'literal': 58, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'literal'}
    instructions[170] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'store'}
    instructions[171] = {5'd0, 4'd8, 4'd0, 16'd108};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'literal': 108, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'literal'}
    instructions[172] = {5'd0, 4'd2, 4'd0, 16'd59};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'literal': 59, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'literal'}
    instructions[173] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'store'}
    instructions[174] = {5'd0, 4'd8, 4'd0, 16'd97};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'literal': 97, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'literal'}
    instructions[175] = {5'd0, 4'd2, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'literal': 60, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'literal'}
    instructions[176] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'store'}
    instructions[177] = {5'd0, 4'd8, 4'd0, 16'd121};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'literal': 121, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'literal'}
    instructions[178] = {5'd0, 4'd2, 4'd0, 16'd61};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'literal': 61, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'literal'}
    instructions[179] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'store'}
    instructions[180] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'literal'}
    instructions[181] = {5'd0, 4'd2, 4'd0, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'literal': 62, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'literal'}
    instructions[182] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'store'}
    instructions[183] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'literal'}
    instructions[184] = {5'd0, 4'd2, 4'd0, 16'd63};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'literal': 63, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'literal'}
    instructions[185] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'store'}
    instructions[186] = {5'd0, 4'd8, 4'd0, 16'd103};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'literal': 103, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'literal'}
    instructions[187] = {5'd0, 4'd2, 4'd0, 16'd64};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'literal': 64, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'literal'}
    instructions[188] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'store'}
    instructions[189] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'literal'}
    instructions[190] = {5'd0, 4'd2, 4'd0, 16'd65};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'literal': 65, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'literal'}
    instructions[191] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'store'}
    instructions[192] = {5'd0, 4'd8, 4'd0, 16'd97};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'literal': 97, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'literal'}
    instructions[193] = {5'd0, 4'd2, 4'd0, 16'd66};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'literal': 66, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'literal'}
    instructions[194] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'store'}
    instructions[195] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'literal'}
    instructions[196] = {5'd0, 4'd2, 4'd0, 16'd67};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'literal': 67, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'literal'}
    instructions[197] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'store'}
    instructions[198] = {5'd0, 4'd8, 4'd0, 16'd100};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'literal': 100, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'literal'}
    instructions[199] = {5'd0, 4'd2, 4'd0, 16'd68};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'literal': 68, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'literal'}
    instructions[200] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'store'}
    instructions[201] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'literal'}
    instructions[202] = {5'd0, 4'd2, 4'd0, 16'd69};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'literal': 69, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'literal'}
    instructions[203] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'store'}
    instructions[204] = {5'd0, 4'd8, 4'd0, 16'd111};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'literal': 111, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'literal'}
    instructions[205] = {5'd0, 4'd2, 4'd0, 16'd70};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'literal': 70, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'literal'}
    instructions[206] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'store'}
    instructions[207] = {5'd0, 4'd8, 4'd0, 16'd58};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'literal': 58, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'literal'}
    instructions[208] = {5'd0, 4'd2, 4'd0, 16'd71};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'literal': 71, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'literal'}
    instructions[209] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'store'}
    instructions[210] = {5'd0, 4'd8, 4'd0, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'literal': 10, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'literal'}
    instructions[211] = {5'd0, 4'd2, 4'd0, 16'd72};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'literal': 72, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'literal'}
    instructions[212] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'store'}
    instructions[213] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'literal'}
    instructions[214] = {5'd0, 4'd2, 4'd0, 16'd73};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'literal': 73, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'literal'}
    instructions[215] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'store'}
    instructions[216] = {5'd0, 4'd8, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 9 {'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 9, 'op': 'literal'}
    instructions[217] = {5'd0, 4'd2, 4'd0, 16'd74};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 9 {'literal': 74, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 9, 'op': 'literal'}
    instructions[218] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 9 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 9, 'op': 'store'}
    instructions[219] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 94 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 94, 'op': 'addl'}
    instructions[220] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 94 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 94, 'op': 'addl'}
    instructions[221] = {5'd3, 4'd6, 4'd0, 16'd223};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 94 {'z': 6, 'label': 223, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 94, 'op': 'call'}
    instructions[222] = {5'd4, 4'd0, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 94 {'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 94, 'op': 'stop'}
    instructions[223] = {5'd1, 4'd3, 4'd3, 16'd76};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 31 {'a': 3, 'literal': 76, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 31, 'op': 'addl'}
    instructions[224] = {5'd0, 4'd8, 4'd0, 16'd58032};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 33 {'literal': 58032, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 33, 'op': 'literal'}
    instructions[225] = {5'd5, 4'd8, 4'd8, 16'd13};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 33 {'a': 8, 'literal': 13, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 33, 'op': 'literal_hi'}
    instructions[226] = {5'd1, 4'd2, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 33 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 33, 'op': 'addl'}
    instructions[227] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 33 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 33, 'op': 'store'}
    instructions[228] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[229] = {5'd1, 4'd2, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 4, 'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'addl'}
    instructions[230] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'store'}
    instructions[231] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[232] = {5'd1, 4'd2, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 4, 'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'addl'}
    instructions[233] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'store'}
    instructions[234] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[235] = {5'd1, 4'd2, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 4, 'literal': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'addl'}
    instructions[236] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'store'}
    instructions[237] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[238] = {5'd1, 4'd2, 4'd4, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 4, 'literal': 4, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'addl'}
    instructions[239] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'store'}
    instructions[240] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[241] = {5'd1, 4'd2, 4'd4, 16'd5};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 4, 'literal': 5, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'addl'}
    instructions[242] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'store'}
    instructions[243] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35, 'op': 'literal'}
    instructions[244] = {5'd1, 4'd2, 4'd4, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35 {'a': 4, 'literal': 6, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35, 'op': 'addl'}
    instructions[245] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35, 'op': 'store'}
    instructions[246] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35, 'op': 'literal'}
    instructions[247] = {5'd1, 4'd2, 4'd4, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35 {'a': 4, 'literal': 7, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35, 'op': 'addl'}
    instructions[248] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35, 'op': 'store'}
    instructions[249] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35, 'op': 'literal'}
    instructions[250] = {5'd1, 4'd2, 4'd4, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35 {'a': 4, 'literal': 8, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35, 'op': 'addl'}
    instructions[251] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35, 'op': 'store'}
    instructions[252] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35, 'op': 'literal'}
    instructions[253] = {5'd1, 4'd2, 4'd4, 16'd9};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35 {'a': 4, 'literal': 9, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35, 'op': 'addl'}
    instructions[254] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35, 'op': 'store'}
    instructions[255] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35, 'op': 'literal'}
    instructions[256] = {5'd1, 4'd2, 4'd4, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35 {'a': 4, 'literal': 10, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35, 'op': 'addl'}
    instructions[257] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35, 'op': 'store'}
    instructions[258] = {5'd0, 4'd8, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[259] = {5'd1, 4'd2, 4'd4, 16'd11};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'a': 4, 'literal': 11, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'addl'}
    instructions[260] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'store'}
    instructions[261] = {5'd0, 4'd8, 4'd0, 16'd57};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'literal': 57, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'literal'}
    instructions[262] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'addl'}
    instructions[263] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'load'}
    instructions[264] = {5'd0, 4'd2, 4'd0, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'literal': 4, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'literal'}
    instructions[265] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'store'}
    instructions[266] = {5'd0, 4'd8, 4'd0, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 39 {'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 39, 'op': 'literal'}
    instructions[267] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 39 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 39, 'op': 'addl'}
    instructions[268] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 39 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 39, 'op': 'load'}
    instructions[269] = {5'd0, 4'd2, 4'd0, 16'd31};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 39 {'literal': 31, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 39, 'op': 'literal'}
    instructions[270] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 39 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 39, 'op': 'store'}
    instructions[271] = {5'd0, 4'd8, 4'd0, 16'd74};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 41 {'literal': 74, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 41, 'op': 'literal'}
    instructions[272] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 41 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 41, 'op': 'addl'}
    instructions[273] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 41 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 41, 'op': 'load'}
    instructions[274] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 41 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 41, 'op': 'store'}
    instructions[275] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 41 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 41, 'op': 'addl'}
    instructions[276] = {5'd0, 4'd8, 4'd0, 16'd16384};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 41 {'literal': 16384, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 41, 'op': 'literal'}
    instructions[277] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 41 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 41, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[278] = {5'd6, 4'd0, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 41 {'a': 3, 'z': 0, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 41, 'op': 'load'}
    instructions[279] = {5'd7, 4'd0, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 41 {'a': 0, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 41, 'op': 'write'}
    instructions[280] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 41 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 41, 'op': 'addl'}
    instructions[281] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'store'}
    instructions[282] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'addl'}
    instructions[283] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'store'}
    instructions[284] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'addl'}
    instructions[285] = {5'd0, 4'd8, 4'd0, 16'd33};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'literal': 33, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'literal'}
    instructions[286] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'store'}
    instructions[287] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'addl'}
    instructions[288] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'addl'}
    instructions[289] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'addl'}
    instructions[290] = {5'd3, 4'd6, 4'd0, 16'd655};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'z': 6, 'label': 655, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'call'}
    instructions[291] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'addl'}
    instructions[292] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[293] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'load'}
    instructions[294] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[295] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'load'}
    instructions[296] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 42, 'op': 'addl'}
    instructions[297] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 43 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 43, 'op': 'store'}
    instructions[298] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 43 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 43, 'op': 'addl'}
    instructions[299] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 43 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 43, 'op': 'store'}
    instructions[300] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 43 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 43, 'op': 'addl'}
    instructions[301] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 43 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 43, 'op': 'addl'}
    instructions[302] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 43 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 43, 'op': 'addl'}
    instructions[303] = {5'd3, 4'd6, 4'd0, 16'd746};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 43 {'z': 6, 'label': 746, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 43, 'op': 'call'}
    instructions[304] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 43 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 43, 'op': 'addl'}
    instructions[305] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 43 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 43, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[306] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 43 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 43, 'op': 'load'}
    instructions[307] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 43 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 43, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[308] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 43 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 43, 'op': 'load'}
    instructions[309] = {5'd0, 4'd2, 4'd0, 16'd5};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 43 {'literal': 5, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 43, 'op': 'literal'}
    instructions[310] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 43 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 43, 'op': 'load'}
    instructions[311] = {5'd1, 4'd2, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 43 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 43, 'op': 'addl'}
    instructions[312] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 43 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 43, 'op': 'store'}
    instructions[313] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'store'}
    instructions[314] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'addl'}
    instructions[315] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'store'}
    instructions[316] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'addl'}
    instructions[317] = {5'd0, 4'd8, 4'd0, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'literal': 7, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'literal'}
    instructions[318] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'store'}
    instructions[319] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'addl'}
    instructions[320] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'addl'}
    instructions[321] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'addl'}
    instructions[322] = {5'd3, 4'd6, 4'd0, 16'd655};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'z': 6, 'label': 655, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'call'}
    instructions[323] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'addl'}
    instructions[324] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[325] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'load'}
    instructions[326] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[327] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'load'}
    instructions[328] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 44, 'op': 'addl'}
    instructions[329] = {5'd0, 4'd8, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45 {'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45, 'op': 'literal'}
    instructions[330] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45, 'op': 'addl'}
    instructions[331] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45, 'op': 'load'}
    instructions[332] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45, 'op': 'store'}
    instructions[333] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45, 'op': 'addl'}
    instructions[334] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45, 'op': 'literal'}
    instructions[335] = {5'd0, 4'd9, 4'd0, 16'd55172};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45 {'literal': 55172, 'z': 9, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45, 'op': 'literal'}
    instructions[336] = {5'd5, 4'd9, 4'd9, 16'd16279};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45 {'a': 9, 'literal': 16279, 'z': 9, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45, 'op': 'literal_hi'}
    instructions[337] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45, 'op': 'store'}
    instructions[338] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45, 'op': 'addl'}
    instructions[339] = {5'd2, 4'd0, 4'd3, 16'd9};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45 {'a': 3, 'comment': 'push', 'b': 9, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45, 'op': 'store'}
    instructions[340] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45, 'op': 'addl'}
    instructions[341] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45, 'op': 'addl'}
    instructions[342] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45, 'op': 'addl'}
    instructions[343] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45, 'op': 'load'}
    instructions[344] = {5'd0, 4'd9, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45 {'literal': 0, 'z': 9, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45, 'op': 'literal'}
    instructions[345] = {5'd8, 4'd9, 4'd9, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45 {'a': 9, 'z': 9, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45, 'op': 'a_hi'}
    instructions[346] = {5'd9, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45 {'a': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45, 'op': 'a_lo'}
    instructions[347] = {5'd10, 4'd0, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45 {'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45, 'op': 'long_to_double'}
    instructions[348] = {5'd9, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45 {'a': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45, 'op': 'a_lo'}
    instructions[349] = {5'd8, 4'd9, 4'd9, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45 {'a': 9, 'z': 9, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45, 'op': 'a_hi'}
    instructions[350] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[351] = {5'd6, 4'd11, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45 {'a': 3, 'z': 11, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45, 'op': 'load'}
    instructions[352] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[353] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45, 'op': 'load'}
    instructions[354] = {5'd11, 4'd11, 4'd11, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45 {'a': 11, 'z': 11, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45, 'op': 'b_hi'}
    instructions[355] = {5'd12, 4'd10, 4'd10, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45 {'a': 10, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45, 'op': 'b_lo'}
    instructions[356] = {5'd8, 4'd9, 4'd9, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45 {'a': 9, 'z': 9, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45, 'op': 'a_hi'}
    instructions[357] = {5'd9, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45 {'a': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45, 'op': 'a_lo'}
    instructions[358] = {5'd13, 4'd0, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45 {'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45, 'op': 'long_float_divide'}
    instructions[359] = {5'd9, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45 {'a': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45, 'op': 'a_lo'}
    instructions[360] = {5'd8, 4'd9, 4'd9, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45 {'a': 9, 'z': 9, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45, 'op': 'a_hi'}
    instructions[361] = {5'd8, 4'd9, 4'd9, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45 {'a': 9, 'z': 9, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45, 'op': 'a_hi'}
    instructions[362] = {5'd9, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45 {'a': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45, 'op': 'a_lo'}
    instructions[363] = {5'd14, 4'd0, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45 {'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45, 'op': 'double_to_long'}
    instructions[364] = {5'd9, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45 {'a': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45, 'op': 'a_lo'}
    instructions[365] = {5'd8, 4'd9, 4'd9, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45 {'a': 9, 'z': 9, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45, 'op': 'a_hi'}
    instructions[366] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[367] = {5'd6, 4'd0, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45 {'a': 3, 'z': 0, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45, 'op': 'load'}
    instructions[368] = {5'd7, 4'd0, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45 {'a': 0, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45, 'op': 'write'}
    instructions[369] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 45, 'op': 'addl'}
    instructions[370] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'store'}
    instructions[371] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'addl'}
    instructions[372] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'store'}
    instructions[373] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'addl'}
    instructions[374] = {5'd0, 4'd8, 4'd0, 16'd58};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'literal': 58, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'literal'}
    instructions[375] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'store'}
    instructions[376] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'addl'}
    instructions[377] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'addl'}
    instructions[378] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'addl'}
    instructions[379] = {5'd3, 4'd6, 4'd0, 16'd655};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'z': 6, 'label': 655, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'call'}
    instructions[380] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'addl'}
    instructions[381] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[382] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'load'}
    instructions[383] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[384] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'load'}
    instructions[385] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'addl'}
    instructions[386] = {5'd1, 4'd8, 4'd4, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 54 {'a': 4, 'literal': 7, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 54, 'op': 'addl'}
    instructions[387] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 54 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 54, 'op': 'addl'}
    instructions[388] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 54 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 54, 'op': 'load'}
    instructions[389] = {5'd1, 4'd2, 4'd4, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 54 {'a': 4, 'literal': 10, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 54, 'op': 'addl'}
    instructions[390] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 54 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 54, 'op': 'store'}
    instructions[391] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 55 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 55, 'op': 'literal'}
    instructions[392] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 55 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 55, 'op': 'addl'}
    instructions[393] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 55 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 55, 'op': 'load'}
    instructions[394] = {5'd15, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 55 {'a': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 55, 'op': 'read'}
    instructions[395] = {5'd1, 4'd2, 4'd4, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 55 {'a': 4, 'literal': 7, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 55, 'op': 'addl'}
    instructions[396] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 55 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 55, 'op': 'store'}
    instructions[397] = {5'd0, 4'd8, 4'd0, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 56 {'literal': 10, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 56, 'op': 'literal'}
    instructions[398] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 56 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 56, 'op': 'store'}
    instructions[399] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 56 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 56, 'op': 'addl'}
    instructions[400] = {5'd1, 4'd8, 4'd4, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 56 {'a': 4, 'literal': 7, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 56, 'op': 'addl'}
    instructions[401] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 56 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 56, 'op': 'addl'}
    instructions[402] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 56 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 56, 'op': 'load'}
    instructions[403] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 56 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 56, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[404] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 56 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 56, 'op': 'load'}
    instructions[405] = {5'd16, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 56 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 56, 'op': 'shift_right'}
    instructions[406] = {5'd1, 4'd2, 4'd4, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 56 {'a': 4, 'literal': 7, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 56, 'op': 'addl'}
    instructions[407] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 56 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 56, 'op': 'store'}
    instructions[408] = {5'd1, 4'd8, 4'd4, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57 {'a': 4, 'literal': 10, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57, 'op': 'addl'}
    instructions[409] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57, 'op': 'addl'}
    instructions[410] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57, 'op': 'load'}
    instructions[411] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57, 'op': 'store'}
    instructions[412] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57, 'op': 'addl'}
    instructions[413] = {5'd1, 4'd8, 4'd4, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57 {'a': 4, 'literal': 7, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57, 'op': 'addl'}
    instructions[414] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57, 'op': 'addl'}
    instructions[415] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57, 'op': 'load'}
    instructions[416] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[417] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57, 'op': 'load'}
    instructions[418] = {5'd17, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57, 'op': 'subtract'}
    instructions[419] = {5'd1, 4'd2, 4'd4, 16'd5};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57 {'a': 4, 'literal': 5, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57, 'op': 'addl'}
    instructions[420] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57, 'op': 'store'}
    instructions[421] = {5'd1, 4'd8, 4'd4, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 60 {'a': 4, 'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 60, 'op': 'addl'}
    instructions[422] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 60 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 60, 'op': 'addl'}
    instructions[423] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 60 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 60, 'op': 'load'}
    instructions[424] = {5'd1, 4'd2, 4'd4, 16'd9};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 60 {'a': 4, 'literal': 9, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 60, 'op': 'addl'}
    instructions[425] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 60 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 60, 'op': 'store'}
    instructions[426] = {5'd1, 4'd8, 4'd4, 16'd5};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 61 {'a': 4, 'literal': 5, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 61, 'op': 'addl'}
    instructions[427] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 61 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 61, 'op': 'addl'}
    instructions[428] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 61 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 61, 'op': 'load'}
    instructions[429] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 61 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 61, 'op': 'store'}
    instructions[430] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 61 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 61, 'op': 'addl'}
    instructions[431] = {5'd0, 4'd8, 4'd0, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 61 {'literal': 10, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 61, 'op': 'literal'}
    instructions[432] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 61 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 61, 'op': 'store'}
    instructions[433] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 61 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 61, 'op': 'addl'}
    instructions[434] = {5'd1, 4'd8, 4'd4, 16'd9};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 61 {'a': 4, 'literal': 9, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 61, 'op': 'addl'}
    instructions[435] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 61 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 61, 'op': 'addl'}
    instructions[436] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 61 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 61, 'op': 'load'}
    instructions[437] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 61 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 61, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[438] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 61 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 61, 'op': 'load'}
    instructions[439] = {5'd16, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 61 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 61, 'op': 'shift_right'}
    instructions[440] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 61 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 61, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[441] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 61 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 61, 'op': 'load'}
    instructions[442] = {5'd18, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 61 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 61, 'op': 'add'}
    instructions[443] = {5'd1, 4'd2, 4'd4, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 61 {'a': 4, 'literal': 6, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 61, 'op': 'addl'}
    instructions[444] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 61 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 61, 'op': 'store'}
    instructions[445] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'addl'}
    instructions[446] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'addl'}
    instructions[447] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'load'}
    instructions[448] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'store'}
    instructions[449] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'addl'}
    instructions[450] = {5'd1, 4'd8, 4'd4, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 4, 'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'addl'}
    instructions[451] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'addl'}
    instructions[452] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'load'}
    instructions[453] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[454] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'load'}
    instructions[455] = {5'd19, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'greater'}
    instructions[456] = {5'd20, 4'd0, 4'd8, 16'd463};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 8, 'label': 463, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'jmp_if_false'}
    instructions[457] = {5'd1, 4'd8, 4'd4, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 4, 'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'addl'}
    instructions[458] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'addl'}
    instructions[459] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'load'}
    instructions[460] = {5'd1, 4'd2, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 4, 'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'addl'}
    instructions[461] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'store'}
    instructions[462] = {5'd21, 4'd0, 4'd0, 16'd463};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'label': 463, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'goto'}
    instructions[463] = {5'd1, 4'd8, 4'd4, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 66 {'a': 4, 'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 66, 'op': 'addl'}
    instructions[464] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 66 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 66, 'op': 'addl'}
    instructions[465] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 66 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 66, 'op': 'load'}
    instructions[466] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 66 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 66, 'op': 'store'}
    instructions[467] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 66 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 66, 'op': 'addl'}
    instructions[468] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 66 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 66, 'op': 'addl'}
    instructions[469] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 66 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 66, 'op': 'addl'}
    instructions[470] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 66 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 66, 'op': 'load'}
    instructions[471] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 66 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 66, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[472] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 66 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 66, 'op': 'load'}
    instructions[473] = {5'd19, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 66 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 66, 'op': 'greater'}
    instructions[474] = {5'd20, 4'd0, 4'd8, 16'd481};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 66 {'a': 8, 'label': 481, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 66, 'op': 'jmp_if_false'}
    instructions[475] = {5'd1, 4'd8, 4'd4, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 66 {'a': 4, 'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 66, 'op': 'addl'}
    instructions[476] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 66 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 66, 'op': 'addl'}
    instructions[477] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 66 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 66, 'op': 'load'}
    instructions[478] = {5'd1, 4'd2, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 66 {'a': 4, 'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 66, 'op': 'addl'}
    instructions[479] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 66 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 66, 'op': 'store'}
    instructions[480] = {5'd21, 4'd0, 4'd0, 16'd481};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 66 {'label': 481, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 66, 'op': 'goto'}
    instructions[481] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 67 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 67, 'op': 'literal'}
    instructions[482] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 67 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 67, 'op': 'store'}
    instructions[483] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 67 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 67, 'op': 'addl'}
    instructions[484] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 67 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 67, 'op': 'addl'}
    instructions[485] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 67 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 67, 'op': 'addl'}
    instructions[486] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 67 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 67, 'op': 'load'}
    instructions[487] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 67 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 67, 'op': 'store'}
    instructions[488] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 67 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 67, 'op': 'addl'}
    instructions[489] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 67 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 67, 'op': 'addl'}
    instructions[490] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 67 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 67, 'op': 'addl'}
    instructions[491] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 67 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 67, 'op': 'load'}
    instructions[492] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 67 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 67, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[493] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 67 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 67, 'op': 'load'}
    instructions[494] = {5'd18, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 67 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 67, 'op': 'add'}
    instructions[495] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 67 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 67, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[496] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 67 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 67, 'op': 'load'}
    instructions[497] = {5'd16, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 67 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 67, 'op': 'shift_right'}
    instructions[498] = {5'd1, 4'd2, 4'd4, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 67 {'a': 4, 'literal': 8, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 67, 'op': 'addl'}
    instructions[499] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 67 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 67, 'op': 'store'}
    instructions[500] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 68 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 68, 'op': 'addl'}
    instructions[501] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 68 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 68, 'op': 'addl'}
    instructions[502] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 68 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 68, 'op': 'load'}
    instructions[503] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 68 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 68, 'op': 'store'}
    instructions[504] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 68 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 68, 'op': 'addl'}
    instructions[505] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 68 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 68, 'op': 'addl'}
    instructions[506] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 68 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 68, 'op': 'addl'}
    instructions[507] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 68 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 68, 'op': 'load'}
    instructions[508] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 68 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 68, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[509] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 68 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 68, 'op': 'load'}
    instructions[510] = {5'd17, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 68 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 68, 'op': 'subtract'}
    instructions[511] = {5'd1, 4'd2, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 68 {'a': 4, 'literal': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 68, 'op': 'addl'}
    instructions[512] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 68 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 68, 'op': 'store'}
    instructions[513] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 69 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 69, 'op': 'literal'}
    instructions[514] = {5'd1, 4'd2, 4'd4, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 69 {'a': 4, 'literal': 4, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 69, 'op': 'addl'}
    instructions[515] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 69 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 69, 'op': 'store'}
    instructions[516] = {5'd0, 4'd8, 4'd0, 16'd256};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 70 {'literal': 256, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 70, 'op': 'literal'}
    instructions[517] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 70 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 70, 'op': 'store'}
    instructions[518] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 70 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 70, 'op': 'addl'}
    instructions[519] = {5'd1, 4'd8, 4'd4, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 70 {'a': 4, 'literal': 4, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 70, 'op': 'addl'}
    instructions[520] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 70 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 70, 'op': 'addl'}
    instructions[521] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 70 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 70, 'op': 'load'}
    instructions[522] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 70 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 70, 'op': 'store'}
    instructions[523] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 70 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 70, 'op': 'addl'}
    instructions[524] = {5'd1, 4'd8, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 70 {'a': 4, 'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 70, 'op': 'addl'}
    instructions[525] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 70 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 70, 'op': 'addl'}
    instructions[526] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 70 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 70, 'op': 'load'}
    instructions[527] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 70 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 70, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[528] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 70 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 70, 'op': 'load'}
    instructions[529] = {5'd16, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 70 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 70, 'op': 'shift_right'}
    instructions[530] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 70 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 70, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[531] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 70 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 70, 'op': 'load'}
    instructions[532] = {5'd19, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 70 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 70, 'op': 'greater'}
    instructions[533] = {5'd20, 4'd0, 4'd8, 16'd553};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73 {'a': 8, 'label': 553, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73, 'op': 'jmp_if_false'}
    instructions[534] = {5'd1, 4'd8, 4'd4, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 71 {'a': 4, 'literal': 4, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 71, 'op': 'addl'}
    instructions[535] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 71 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 71, 'op': 'addl'}
    instructions[536] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 71 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 71, 'op': 'load'}
    instructions[537] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 71 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 71, 'op': 'store'}
    instructions[538] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 71 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 71, 'op': 'addl'}
    instructions[539] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 71 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 71, 'op': 'literal'}
    instructions[540] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 71 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 71, 'op': 'store'}
    instructions[541] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 71 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 71, 'op': 'addl'}
    instructions[542] = {5'd1, 4'd8, 4'd4, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 71 {'a': 4, 'literal': 4, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 71, 'op': 'addl'}
    instructions[543] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 71 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 71, 'op': 'addl'}
    instructions[544] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 71 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 71, 'op': 'load'}
    instructions[545] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 71 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 71, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[546] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 71 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 71, 'op': 'load'}
    instructions[547] = {5'd18, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 71 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 71, 'op': 'add'}
    instructions[548] = {5'd1, 4'd2, 4'd4, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 71 {'a': 4, 'literal': 4, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 71, 'op': 'addl'}
    instructions[549] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 71 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 71, 'op': 'store'}
    instructions[550] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 71 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 71, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[551] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 71 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 71, 'op': 'load'}
    instructions[552] = {5'd21, 4'd0, 4'd0, 16'd554};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73 {'label': 554, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73, 'op': 'goto'}
    instructions[553] = {5'd21, 4'd0, 4'd0, 16'd555};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73 {'label': 555, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73, 'op': 'goto'}
    instructions[554] = {5'd21, 4'd0, 4'd0, 16'd516};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 70 {'label': 516, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 70, 'op': 'goto'}
    instructions[555] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73, 'op': 'store'}
    instructions[556] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73, 'op': 'addl'}
    instructions[557] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73, 'op': 'store'}
    instructions[558] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73, 'op': 'addl'}
    instructions[559] = {5'd1, 4'd8, 4'd4, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73 {'a': 4, 'literal': 4, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73, 'op': 'addl'}
    instructions[560] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73, 'op': 'addl'}
    instructions[561] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73, 'op': 'load'}
    instructions[562] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73, 'op': 'store'}
    instructions[563] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73, 'op': 'addl'}
    instructions[564] = {5'd1, 4'd8, 4'd4, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73 {'a': 4, 'literal': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73, 'op': 'addl'}
    instructions[565] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73, 'op': 'addl'}
    instructions[566] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73, 'op': 'load'}
    instructions[567] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73, 'op': 'store'}
    instructions[568] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73, 'op': 'addl'}
    instructions[569] = {5'd1, 4'd8, 4'd4, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73 {'a': 4, 'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73, 'op': 'addl'}
    instructions[570] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73, 'op': 'addl'}
    instructions[571] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73, 'op': 'load'}
    instructions[572] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[573] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73, 'op': 'load'}
    instructions[574] = {5'd17, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73, 'op': 'subtract'}
    instructions[575] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[576] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73, 'op': 'load'}
    instructions[577] = {5'd16, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73, 'op': 'shift_right'}
    instructions[578] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73, 'op': 'store'}
    instructions[579] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73, 'op': 'addl'}
    instructions[580] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73, 'op': 'addl'}
    instructions[581] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73, 'op': 'addl'}
    instructions[582] = {5'd3, 4'd6, 4'd0, 16'd873};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73 {'z': 6, 'label': 873, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73, 'op': 'call'}
    instructions[583] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73, 'op': 'addl'}
    instructions[584] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[585] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73, 'op': 'load'}
    instructions[586] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[587] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73, 'op': 'load'}
    instructions[588] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 73, 'op': 'addl'}
    instructions[589] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74, 'op': 'literal'}
    instructions[590] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74, 'op': 'store'}
    instructions[591] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74, 'op': 'addl'}
    instructions[592] = {5'd1, 4'd8, 4'd4, 16'd11};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74 {'a': 4, 'literal': 11, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74, 'op': 'addl'}
    instructions[593] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74, 'op': 'addl'}
    instructions[594] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74, 'op': 'load'}
    instructions[595] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74, 'op': 'store'}
    instructions[596] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74, 'op': 'addl'}
    instructions[597] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74, 'op': 'literal'}
    instructions[598] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74, 'op': 'store'}
    instructions[599] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74, 'op': 'addl'}
    instructions[600] = {5'd1, 4'd8, 4'd4, 16'd11};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74 {'a': 4, 'literal': 11, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74, 'op': 'addl'}
    instructions[601] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74, 'op': 'addl'}
    instructions[602] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74, 'op': 'load'}
    instructions[603] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[604] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74, 'op': 'load'}
    instructions[605] = {5'd17, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74, 'op': 'subtract'}
    instructions[606] = {5'd1, 4'd2, 4'd4, 16'd11};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74 {'a': 4, 'literal': 11, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74, 'op': 'addl'}
    instructions[607] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74, 'op': 'store'}
    instructions[608] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[609] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74, 'op': 'load'}
    instructions[610] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[611] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74, 'op': 'load'}
    instructions[612] = {5'd22, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74, 'op': 'equal'}
    instructions[613] = {5'd20, 4'd0, 4'd8, 16'd651};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74 {'a': 8, 'label': 651, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74, 'op': 'jmp_if_false'}
    instructions[614] = {5'd0, 4'd8, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 75 {'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 75, 'op': 'literal'}
    instructions[615] = {5'd1, 4'd2, 4'd4, 16'd11};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 75 {'a': 4, 'literal': 11, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 75, 'op': 'addl'}
    instructions[616] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 75 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 75, 'op': 'store'}
    instructions[617] = {5'd0, 4'd8, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 76 {'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 76, 'op': 'literal'}
    instructions[618] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 76 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 76, 'op': 'store'}
    instructions[619] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 76 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 76, 'op': 'addl'}
    instructions[620] = {5'd1, 4'd8, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 76 {'a': 4, 'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 76, 'op': 'addl'}
    instructions[621] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 76 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 76, 'op': 'addl'}
    instructions[622] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 76 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 76, 'op': 'load'}
    instructions[623] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 76 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 76, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[624] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 76 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 76, 'op': 'load'}
    instructions[625] = {5'd19, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 76 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 76, 'op': 'greater'}
    instructions[626] = {5'd20, 4'd0, 4'd8, 16'd650};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 76 {'a': 8, 'label': 650, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 76, 'op': 'jmp_if_false'}
    instructions[627] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 77 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 77, 'op': 'literal'}
    instructions[628] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 77 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 77, 'op': 'store'}
    instructions[629] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 77 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 77, 'op': 'addl'}
    instructions[630] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 77 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 77, 'op': 'addl'}
    instructions[631] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 77 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 77, 'op': 'addl'}
    instructions[632] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 77 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 77, 'op': 'load'}
    instructions[633] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 77 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 77, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[634] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 77 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 77, 'op': 'load'}
    instructions[635] = {5'd17, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 77 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 77, 'op': 'subtract'}
    instructions[636] = {5'd1, 4'd2, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 77 {'a': 4, 'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 77, 'op': 'addl'}
    instructions[637] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 77 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 77, 'op': 'store'}
    instructions[638] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 78 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 78, 'op': 'literal'}
    instructions[639] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 78 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 78, 'op': 'store'}
    instructions[640] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 78 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 78, 'op': 'addl'}
    instructions[641] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 78 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 78, 'op': 'addl'}
    instructions[642] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 78 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 78, 'op': 'addl'}
    instructions[643] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 78 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 78, 'op': 'load'}
    instructions[644] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 78 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 78, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[645] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 78 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 78, 'op': 'load'}
    instructions[646] = {5'd18, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 78 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 78, 'op': 'add'}
    instructions[647] = {5'd1, 4'd2, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 78 {'a': 4, 'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 78, 'op': 'addl'}
    instructions[648] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 78 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 78, 'op': 'store'}
    instructions[649] = {5'd21, 4'd0, 4'd0, 16'd650};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 76 {'label': 650, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 76, 'op': 'goto'}
    instructions[650] = {5'd21, 4'd0, 4'd0, 16'd651};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74 {'label': 651, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 74, 'op': 'goto'}
    instructions[651] = {5'd21, 4'd0, 4'd0, 16'd386};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 48 {'label': 386, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 48, 'op': 'goto'}
    instructions[652] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 31 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 31, 'op': 'addl'}
    instructions[653] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 31 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 31, 'op': 'addl'}
    instructions[654] = {5'd23, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 31 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 31, 'op': 'return'}
    instructions[655] = {5'd1, 4'd3, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73 {'a': 3, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73, 'op': 'addl'}
    instructions[656] = {5'd2, 4'd0, 4'd3, 16'd6};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'store'}
    instructions[657] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[658] = {5'd2, 4'd0, 4'd3, 16'd7};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'store'}
    instructions[659] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[660] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[661] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[662] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'load'}
    instructions[663] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'store'}
    instructions[664] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[665] = {5'd0, 4'd8, 4'd0, 16'd4};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'literal': 4, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'literal'}
    instructions[666] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[667] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'load'}
    instructions[668] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'store'}
    instructions[669] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[670] = {5'd1, 4'd7, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 4, 'literal': 0, 'z': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[671] = {5'd1, 4'd4, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[672] = {5'd3, 4'd6, 4'd0, 16'd682};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'z': 6, 'label': 682, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'call'}
    instructions[673] = {5'd1, 4'd3, 4'd3, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': -2, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[674] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[675] = {5'd6, 4'd7, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'z': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'load'}
    instructions[676] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[677] = {5'd6, 4'd6, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'z': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'load'}
    instructions[678] = {5'd1, 4'd3, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[679] = {5'd1, 4'd3, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73 {'a': 4, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73, 'op': 'addl'}
    instructions[680] = {5'd1, 4'd4, 4'd7, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73 {'a': 7, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73, 'op': 'addl'}
    instructions[681] = {5'd23, 4'd0, 4'd6, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73 {'a': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73, 'op': 'return'}
    instructions[682] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23, 'op': 'addl'}
    instructions[683] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 24 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 24, 'op': 'literal'}
    instructions[684] = {5'd1, 4'd2, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 24 {'a': 4, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 24, 'op': 'addl'}
    instructions[685] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 24 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 24, 'op': 'store'}
    instructions[686] = {5'd1, 4'd8, 4'd4, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 4, 'literal': -2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'addl'}
    instructions[687] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'addl'}
    instructions[688] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'load'}
    instructions[689] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'store'}
    instructions[690] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'addl'}
    instructions[691] = {5'd1, 4'd8, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 4, 'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'addl'}
    instructions[692] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'addl'}
    instructions[693] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'load'}
    instructions[694] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[695] = {5'd6, 4'd2, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 3, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'load'}
    instructions[696] = {5'd18, 4'd8, 4'd8, 16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 8, 'z': 8, 'b': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'add'}
    instructions[697] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'addl'}
    instructions[698] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'load'}
    instructions[699] = {5'd20, 4'd0, 4'd8, 16'd741};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 29 {'a': 8, 'label': 741, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 29, 'op': 'jmp_if_false'}
    instructions[700] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[701] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[702] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'load'}
    instructions[703] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'store'}
    instructions[704] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[705] = {5'd1, 4'd8, 4'd4, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 4, 'literal': -2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[706] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[707] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'load'}
    instructions[708] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'store'}
    instructions[709] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[710] = {5'd1, 4'd8, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 4, 'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[711] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[712] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'load'}
    instructions[713] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[714] = {5'd6, 4'd2, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'load'}
    instructions[715] = {5'd18, 4'd8, 4'd8, 16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 8, 'z': 8, 'b': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'add'}
    instructions[716] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[717] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'load'}
    instructions[718] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[719] = {5'd6, 4'd0, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'z': 0, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'load'}
    instructions[720] = {5'd7, 4'd0, 4'd0, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 0, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'write'}
    instructions[721] = {5'd1, 4'd3, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[722] = {5'd1, 4'd8, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 4, 'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[723] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[724] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'load'}
    instructions[725] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'store'}
    instructions[726] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[727] = {5'd0, 4'd8, 4'd0, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'literal': 1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'literal'}
    instructions[728] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'store'}
    instructions[729] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[730] = {5'd1, 4'd8, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 4, 'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[731] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[732] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'load'}
    instructions[733] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[734] = {5'd6, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'load'}
    instructions[735] = {5'd18, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'add'}
    instructions[736] = {5'd1, 4'd2, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 4, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[737] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'store'}
    instructions[738] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[739] = {5'd6, 4'd8, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'load'}
    instructions[740] = {5'd21, 4'd0, 4'd0, 16'd742};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 29 {'label': 742, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 29, 'op': 'goto'}
    instructions[741] = {5'd21, 4'd0, 4'd0, 16'd743};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 29 {'label': 743, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 29, 'op': 'goto'}
    instructions[742] = {5'd21, 4'd0, 4'd0, 16'd686};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'label': 686, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'goto'}
    instructions[743] = {5'd1, 4'd3, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23 {'a': 4, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23, 'op': 'addl'}
    instructions[744] = {5'd1, 4'd4, 4'd7, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23 {'a': 7, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23, 'op': 'addl'}
    instructions[745] = {5'd23, 4'd0, 4'd6, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23 {'a': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23, 'op': 'return'}
    instructions[746] = {5'd1, 4'd3, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 155 {'a': 3, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 155, 'op': 'addl'}
    instructions[747] = {5'd2, 4'd0, 4'd3, 16'd6};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'op': 'store'}
    instructions[748] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'op': 'addl'}
    instructions[749] = {5'd2, 4'd0, 4'd3, 16'd7};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'op': 'store'}
    instructions[750] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'op': 'addl'}
    instructions[751] = {5'd0, 4'd8, 4'd0, 16'd31};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'literal': 31, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'op': 'literal'}
    instructions[752] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'op': 'addl'}
    instructions[753] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'op': 'load'}
    instructions[754] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'op': 'store'}
    instructions[755] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'op': 'addl'}
    instructions[756] = {5'd1, 4'd7, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'a': 4, 'literal': 0, 'z': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'op': 'addl'}
    instructions[757] = {5'd1, 4'd4, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'a': 3, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'op': 'addl'}
    instructions[758] = {5'd3, 4'd6, 4'd0, 16'd771};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'z': 6, 'label': 771, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'op': 'call'}
    instructions[759] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'a': 3, 'literal': -1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'op': 'addl'}
    instructions[760] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[761] = {5'd6, 4'd7, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'a': 3, 'z': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'op': 'load'}
    instructions[762] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[763] = {5'd6, 4'd6, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'a': 3, 'z': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'op': 'load'}
    instructions[764] = {5'd0, 4'd2, 4'd0, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'literal': 1, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'op': 'literal'}
    instructions[765] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'op': 'load'}
    instructions[766] = {5'd0, 4'd2, 4'd0, 16'd5};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'literal': 5, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'op': 'literal'}
    instructions[767] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'op': 'store'}
    instructions[768] = {5'd1, 4'd3, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'a': 4, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'op': 'addl'}
    instructions[769] = {5'd1, 4'd4, 4'd7, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'a': 7, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'op': 'addl'}
    instructions[770] = {5'd23, 4'd0, 4'd6, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'a': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'op': 'return'}
    instructions[771] = {5'd1, 4'd3, 4'd3, 16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 26 {'a': 3, 'literal': 2, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 26, 'op': 'addl'}
    instructions[772] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 29 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 29, 'op': 'literal'}
    instructions[773] = {5'd1, 4'd2, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 29 {'a': 4, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 29, 'op': 'addl'}
    instructions[774] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 29 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 29, 'op': 'store'}
    instructions[775] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 31 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 31, 'op': 'addl'}
    instructions[776] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 31 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 31, 'op': 'addl'}
    instructions[777] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 31 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 31, 'op': 'load'}
    instructions[778] = {5'd15, 4'd8, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 31 {'a': 8, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 31, 'op': 'read'}
    instructions[779] = {5'd1, 4'd2, 4'd4, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 31 {'a': 4, 'literal': 1, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 31, 'op': 'addl'}
    instructions[780] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 31 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 31, 'op': 'store'}
    instructions[781] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'literal'}
    instructions[782] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'store'}
    instructions[783] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'addl'}
    instructions[784] = {5'd2, 4'd0, 4'd3, 16'd6};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'store'}
    instructions[785] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'addl'}
    instructions[786] = {5'd2, 4'd0, 4'd3, 16'd7};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'store'}
    instructions[787] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'addl'}
    instructions[788] = {5'd1, 4'd8, 4'd4, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'a': 4, 'literal': 1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'addl'}
    instructions[789] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'addl'}
    instructions[790] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'load'}
    instructions[791] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'store'}
    instructions[792] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'addl'}
    instructions[793] = {5'd1, 4'd7, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'a': 4, 'literal': 0, 'z': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'addl'}
    instructions[794] = {5'd1, 4'd4, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'a': 3, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'addl'}
    instructions[795] = {5'd3, 4'd6, 4'd0, 16'd848};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'z': 6, 'label': 848, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'call'}
    instructions[796] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'a': 3, 'literal': -1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'addl'}
    instructions[797] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[798] = {5'd6, 4'd7, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'a': 3, 'z': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'load'}
    instructions[799] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[800] = {5'd6, 4'd6, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'a': 3, 'z': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'load'}
    instructions[801] = {5'd0, 4'd2, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'literal'}
    instructions[802] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'load'}
    instructions[803] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[804] = {5'd6, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'load'}
    instructions[805] = {5'd22, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'equal'}
    instructions[806] = {5'd20, 4'd0, 4'd8, 16'd809};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'a': 8, 'label': 809, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'jmp_if_false'}
    instructions[807] = {5'd21, 4'd0, 4'd0, 16'd840};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'label': 840, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'goto'}
    instructions[808] = {5'd21, 4'd0, 4'd0, 16'd809};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'label': 809, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'goto'}
    instructions[809] = {5'd0, 4'd8, 4'd0, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 33 {'literal': 10, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 33, 'op': 'literal'}
    instructions[810] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 33 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 33, 'op': 'store'}
    instructions[811] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 33 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 33, 'op': 'addl'}
    instructions[812] = {5'd1, 4'd8, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 33 {'a': 4, 'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 33, 'op': 'addl'}
    instructions[813] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 33 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 33, 'op': 'addl'}
    instructions[814] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 33 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 33, 'op': 'load'}
    instructions[815] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 33 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 33, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[816] = {5'd6, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 33 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 33, 'op': 'load'}
    instructions[817] = {5'd24, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 33 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 33, 'op': 'multiply'}
    instructions[818] = {5'd1, 4'd2, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 33 {'a': 4, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 33, 'op': 'addl'}
    instructions[819] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 33 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 33, 'op': 'store'}
    instructions[820] = {5'd0, 4'd8, 4'd0, 16'd48};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34 {'literal': 48, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34, 'op': 'literal'}
    instructions[821] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34, 'op': 'store'}
    instructions[822] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34, 'op': 'addl'}
    instructions[823] = {5'd1, 4'd8, 4'd4, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34 {'a': 4, 'literal': 1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34, 'op': 'addl'}
    instructions[824] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34, 'op': 'addl'}
    instructions[825] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34, 'op': 'load'}
    instructions[826] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[827] = {5'd6, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34, 'op': 'load'}
    instructions[828] = {5'd17, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34, 'op': 'subtract'}
    instructions[829] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34, 'op': 'store'}
    instructions[830] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34, 'op': 'addl'}
    instructions[831] = {5'd1, 4'd8, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34 {'a': 4, 'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34, 'op': 'addl'}
    instructions[832] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34, 'op': 'addl'}
    instructions[833] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34, 'op': 'load'}
    instructions[834] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[835] = {5'd6, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34, 'op': 'load'}
    instructions[836] = {5'd18, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34, 'op': 'add'}
    instructions[837] = {5'd1, 4'd2, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34 {'a': 4, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34, 'op': 'addl'}
    instructions[838] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34, 'op': 'store'}
    instructions[839] = {5'd21, 4'd0, 4'd0, 16'd775};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 30 {'label': 775, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 30, 'op': 'goto'}
    instructions[840] = {5'd1, 4'd8, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 36 {'a': 4, 'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 36, 'op': 'addl'}
    instructions[841] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 36 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 36, 'op': 'addl'}
    instructions[842] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 36 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 36, 'op': 'load'}
    instructions[843] = {5'd0, 4'd2, 4'd0, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 36 {'literal': 1, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 36, 'op': 'literal'}
    instructions[844] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 36 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 36, 'op': 'store'}
    instructions[845] = {5'd1, 4'd3, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 36 {'a': 4, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 36, 'op': 'addl'}
    instructions[846] = {5'd1, 4'd4, 4'd7, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 36 {'a': 7, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 36, 'op': 'addl'}
    instructions[847] = {5'd23, 4'd0, 4'd6, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 36 {'a': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 36, 'op': 'return'}
    instructions[848] = {5'd1, 4'd3, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 86 {'a': 3, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 86, 'op': 'addl'}
    instructions[849] = {5'd0, 4'd8, 4'd0, 16'd48};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'literal': 48, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'op': 'literal'}
    instructions[850] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'op': 'store'}
    instructions[851] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'op': 'addl'}
    instructions[852] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'op': 'addl'}
    instructions[853] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'op': 'addl'}
    instructions[854] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'op': 'load'}
    instructions[855] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[856] = {5'd6, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'op': 'load'}
    instructions[857] = {5'd25, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'op': 'greater_equal'}
    instructions[858] = {5'd20, 4'd0, 4'd8, 16'd868};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'a': 8, 'label': 868, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'op': 'jmp_if_false'}
    instructions[859] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'op': 'addl'}
    instructions[860] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'op': 'addl'}
    instructions[861] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'op': 'load'}
    instructions[862] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'op': 'store'}
    instructions[863] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'op': 'addl'}
    instructions[864] = {5'd0, 4'd8, 4'd0, 16'd57};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'literal': 57, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'op': 'literal'}
    instructions[865] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[866] = {5'd6, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'op': 'load'}
    instructions[867] = {5'd25, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'op': 'greater_equal'}
    instructions[868] = {5'd0, 4'd2, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'op': 'literal'}
    instructions[869] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'op': 'store'}
    instructions[870] = {5'd1, 4'd3, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'a': 4, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'op': 'addl'}
    instructions[871] = {5'd1, 4'd4, 4'd7, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'a': 7, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'op': 'addl'}
    instructions[872] = {5'd23, 4'd0, 4'd6, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'a': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'op': 'return'}
    instructions[873] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 25 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 25, 'op': 'addl'}
    instructions[874] = {5'd0, 4'd8, 4'd0, 16'd127};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 26 {'literal': 127, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 26, 'op': 'literal'}
    instructions[875] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 26 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 26, 'op': 'store'}
    instructions[876] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 26 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 26, 'op': 'addl'}
    instructions[877] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 26 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 26, 'op': 'addl'}
    instructions[878] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 26 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 26, 'op': 'addl'}
    instructions[879] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 26 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 26, 'op': 'load'}
    instructions[880] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 26 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 26, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[881] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 26 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 26, 'op': 'load'}
    instructions[882] = {5'd19, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 26 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 26, 'op': 'greater'}
    instructions[883] = {5'd20, 4'd0, 4'd8, 16'd888};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 26 {'a': 8, 'label': 888, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 26, 'op': 'jmp_if_false'}
    instructions[884] = {5'd0, 4'd8, 4'd0, 16'd127};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 26 {'literal': 127, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 26, 'op': 'literal'}
    instructions[885] = {5'd1, 4'd2, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 26 {'a': 4, 'literal': -1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 26, 'op': 'addl'}
    instructions[886] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 26 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 26, 'op': 'store'}
    instructions[887] = {5'd21, 4'd0, 4'd0, 16'd888};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 26 {'label': 888, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 26, 'op': 'goto'}
    instructions[888] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27, 'op': 'addl'}
    instructions[889] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27, 'op': 'addl'}
    instructions[890] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27, 'op': 'load'}
    instructions[891] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27, 'op': 'store'}
    instructions[892] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27, 'op': 'addl'}
    instructions[893] = {5'd0, 4'd8, 4'd0, 16'd65408};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27 {'literal': 65408, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27, 'op': 'literal'}
    instructions[894] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[895] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27, 'op': 'load'}
    instructions[896] = {5'd19, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27, 'op': 'greater'}
    instructions[897] = {5'd20, 4'd0, 4'd8, 16'd902};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27 {'a': 8, 'label': 902, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27, 'op': 'jmp_if_false'}
    instructions[898] = {5'd0, 4'd8, 4'd0, 16'd65408};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27 {'literal': 65408, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27, 'op': 'literal'}
    instructions[899] = {5'd1, 4'd2, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27 {'a': 4, 'literal': -1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27, 'op': 'addl'}
    instructions[900] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27, 'op': 'store'}
    instructions[901] = {5'd21, 4'd0, 4'd0, 16'd902};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27 {'label': 902, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27, 'op': 'goto'}
    instructions[902] = {5'd0, 4'd8, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28 {'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28, 'op': 'literal'}
    instructions[903] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28, 'op': 'addl'}
    instructions[904] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28, 'op': 'load'}
    instructions[905] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28, 'op': 'store'}
    instructions[906] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28, 'op': 'addl'}
    instructions[907] = {5'd0, 4'd8, 4'd0, 16'd128};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28 {'literal': 128, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28, 'op': 'literal'}
    instructions[908] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28, 'op': 'store'}
    instructions[909] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28, 'op': 'addl'}
    instructions[910] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28, 'op': 'addl'}
    instructions[911] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28, 'op': 'addl'}
    instructions[912] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28, 'op': 'load'}
    instructions[913] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[914] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28, 'op': 'load'}
    instructions[915] = {5'd18, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28, 'op': 'add'}
    instructions[916] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[917] = {5'd6, 4'd0, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28 {'a': 3, 'z': 0, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28, 'op': 'load'}
    instructions[918] = {5'd7, 4'd0, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28 {'a': 0, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28, 'op': 'write'}
    instructions[919] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28, 'op': 'addl'}
    instructions[920] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 25 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 25, 'op': 'addl'}
    instructions[921] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 25 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 25, 'op': 'addl'}
    instructions[922] = {5'd23, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 25 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 25, 'op': 'return'}
  end

  
  always @(posedge clk)
  begin
    load_data <= memory[load_address];
    if(store_enable && state == execute) begin
      memory[store_address] <= store_data;
    end
  end


  //////////////////////////////////////////////////////////////////////////////
  // PIPELINE STAGE 1 -- FETCH INSTRUCTION
  //                                                                            
  
  always @(posedge clk)
  begin
    //implement memory for instructions
    if (state == instruction_fetch || state == operand_fetch || state == execute) begin
      instruction <= instructions[program_counter];
      program_counter_1 <= program_counter;
    end
  end

  assign opcode    = instruction[28:24];
  assign address_z = instruction[23:20];
  assign address_a = instruction[19:16];
  assign address_b = instruction[3:0];
  assign literal   = instruction[15:0];

  //////////////////////////////////////////////////////////////////////////////
  // PIPELINE STAGE 2 -- FETCH OPERANDS
  //                                                                            
  
  always @(posedge clk)
  begin
    if (write_enable) begin
      registers[address_z_3] <= result;
    end
    if (state == operand_fetch || state == execute) begin
      opcode_2 <= opcode;
      literal_2 <= literal;
      address_a_2 <= address_a;
      address_b_2 <= address_b;
      address_z_2 <= address_z;
      program_counter_2 <= program_counter_1;
    end
  end
  assign register_a = registers[address_a_2];
  assign register_b = registers[address_b_2];
  assign operand_a = (address_a_2 == address_z_3 && write_enable)?result:register_a;
  assign operand_b = (address_b_2 == address_z_3 && write_enable)?result:register_b;
  assign store_address = operand_a;
  assign load_address = operand_a;
  assign store_data = operand_b;
  assign store_enable = (opcode_2==2);

  //////////////////////////////////////////////////////////////////////////////
  // PIPELINE STAGE 3 -- EXECUTE
  //                                                                            
  
  always @(posedge clk)
  begin

  write_enable <= 0;
  timer_clock <= timer_clock + 1;
  case(state)

    //instruction_fetch
    instruction_fetch: begin
      program_counter <= program_counter + 1;
      state <= operand_fetch;
    end
    //operand_fetch
    operand_fetch: begin
      program_counter <= program_counter + 1;
      state <= execute;
    end
    //execute
    execute: begin
      program_counter <= program_counter + 1;
      address_z_3 <= address_z_2;
      case(opcode_2)

        //literal
        16'd0:
        begin
          result<=$signed(literal_2);
          write_enable <= 1;
        end

        //addl
        16'd1:
        begin
          result<=operand_a + literal_2;
          write_enable <= 1;
        end

        //store
        16'd2:
        begin
        end

        //call
        16'd3:
        begin
          result <= program_counter_2 + 1;
          write_enable <= 1;
          program_counter <= literal_2;
          state <= instruction_fetch;
        end

        //stop
        16'd4:
        begin
        state <= stop;
        end

        //literal_hi
        16'd5:
        begin
          result<= {literal_2, operand_a[15:0]};
          write_enable <= 1;
        end

        //load
        16'd6:
        begin
          state <= load;
        end

        //write
        16'd7:
        begin
          state <= write;
          write_output <= operand_a;
          write_value <= operand_b;
        end

        //a_hi
        16'd8:
        begin
          a_hi <= operand_a;
          result <= a_hi;
          write_enable <= 1;
        end

        //a_lo
        16'd9:
        begin
          a_lo <= operand_a;
          result <= a_lo;
          write_enable <= 1;
        end

        //long_to_double
        16'd10:
        begin
          long_to_double_in <= {a_hi, a_lo};
          state <= long_to_double_write_a;
        end

        //b_hi
        16'd11:
        begin
          b_hi <= operand_a;
          result <= b_hi;
          write_enable <= 1;
        end

        //b_lo
        16'd12:
        begin
          b_lo <= operand_a;
          result <= b_lo;
          write_enable <= 1;
        end

        //long_float_divide
        16'd13:
        begin
          double_divider_a <= {a_hi, a_lo};
          double_divider_b <= {b_hi, b_lo};
          state <= double_divider_write_a;
        end

        //double_to_long
        16'd14:
        begin
          double_to_long_in <= {a_hi, a_lo};
          state <= double_to_long_write_a;
        end

        //read
        16'd15:
        begin
          state <= read;
          read_input <= operand_a;
        end

        //shift_right
        16'd16:
        begin
          if(operand_b < 32) begin
            result <= $signed(operand_a) >>> operand_b;
            carry <= operand_a << (32-operand_b);
          end else begin
            result <= operand_a[31]?-1:0;
            carry <= operand_a;
          end
          write_enable <= 1;
        end

        //subtract
        16'd17:
        begin
          long_result = operand_a + (~operand_b) + 1;
          result <= long_result[31:0];
          carry[0] <= ~long_result[32];
          write_enable <= 1;
        end

        //add
        16'd18:
        begin
          long_result = operand_a + operand_b;
          result <= long_result[31:0];
          carry[0] <= long_result[32];
          write_enable <= 1;
        end

        //greater
        16'd19:
        begin
          result <= $signed(operand_a) > $signed(operand_b);
          write_enable <= 1;
        end

        //jmp_if_false
        16'd20:
        begin
          if (operand_a == 0) begin
            program_counter <= literal_2;
            state <= instruction_fetch;
          end
        end

        //goto
        16'd21:
        begin
          program_counter <= literal_2;
          state <= instruction_fetch;
        end

        //equal
        16'd22:
        begin
          result <= operand_a == operand_b;
          write_enable <= 1;
        end

        //return
        16'd23:
        begin
          program_counter <= operand_a;
          state <= instruction_fetch;
        end

        //multiply
        16'd24:
        begin
          product_a <= operand_a[15:0]  * operand_b[15:0];
          product_b <= operand_a[15:0]  * operand_b[31:16];
          product_c <= operand_a[31:16] * operand_b[15:0];
          product_d <= operand_a[31:16] * operand_b[31:16];
          state <= multiply;
        end

        //greater_equal
        16'd25:
        begin
          result <= $signed(operand_a) >= $signed(operand_b);
          write_enable <= 1;
        end

      endcase

    end

    multiply:
    begin
      long_result = product_a +
                    (product_b << 16) +
                    (product_c << 16) +
                    (product_d << 32);
      result <= long_result[31:0];
      carry <= long_result[63:32];
      write_enable <= 1;
      state <= execute;
    end

    read:
    begin
      case(read_input)
      0:
      begin
        s_input_eth_in_ack <= 1;
        if (s_input_eth_in_ack && input_eth_in_stb) begin
          result <= input_eth_in;
          write_enable <= 1;
          s_input_eth_in_ack <= 0;
          state <= execute;
        end
      end
      1:
      begin
        s_input_audio_in_ack <= 1;
        if (s_input_audio_in_ack && input_audio_in_stb) begin
          result <= input_audio_in;
          write_enable <= 1;
          s_input_audio_in_ack <= 0;
          state <= execute;
        end
      end
      2:
      begin
        s_input_rs232_rx_ack <= 1;
        if (s_input_rs232_rx_ack && input_rs232_rx_stb) begin
          result <= input_rs232_rx;
          write_enable <= 1;
          s_input_rs232_rx_ack <= 0;
          state <= execute;
        end
      end
      endcase
    end

    write:
    begin
      case(write_output)
      3:
      begin
        s_output_eth_out_stb <= 1;
        s_output_eth_out <= write_value;
        if (output_eth_out_ack && s_output_eth_out_stb) begin
          s_output_eth_out_stb <= 0;
          state <= execute;
        end
      end
      4:
      begin
        s_output_audio_out_stb <= 1;
        s_output_audio_out <= write_value;
        if (output_audio_out_ack && s_output_audio_out_stb) begin
          s_output_audio_out_stb <= 0;
          state <= execute;
        end
      end
      5:
      begin
        s_output_frequency_out_stb <= 1;
        s_output_frequency_out <= write_value;
        if (output_frequency_out_ack && s_output_frequency_out_stb) begin
          s_output_frequency_out_stb <= 0;
          state <= execute;
        end
      end
      6:
      begin
        s_output_samples_out_stb <= 1;
        s_output_samples_out <= write_value;
        if (output_samples_out_ack && s_output_samples_out_stb) begin
          s_output_samples_out_stb <= 0;
          state <= execute;
        end
      end
      7:
      begin
        s_output_rs232_tx_stb <= 1;
        s_output_rs232_tx <= write_value;
        if (output_rs232_tx_ack && s_output_rs232_tx_stb) begin
          s_output_rs232_tx_stb <= 0;
          state <= execute;
        end
      end
      endcase
    end

    load:
    begin
        result <= load_data;
        write_enable <= 1;
        state <= execute;
    end

    wait_state:
    begin
      if (timer) begin
        timer <= timer - 1;
      end else begin
        state <= execute;
      end
    end

    stop:
    begin
    end

    double_divider_write_a:
    begin
      double_divider_a_stb <= 1;
      if (double_divider_a_stb && double_divider_a_ack) begin
        double_divider_a_stb <= 0;
        state <= double_divider_write_b;
      end
    end

    double_divider_write_b:
    begin
      double_divider_b_stb <= 1;
      if (double_divider_b_stb && double_divider_b_ack) begin
        double_divider_b_stb <= 0;
        state <= double_divider_read_z;
      end
    end

    double_divider_read_z:
    begin
      double_divider_z_ack <= 1;
      if (double_divider_z_stb && double_divider_z_ack) begin
        a_lo <= double_divider_z[31:0];
        a_hi <= double_divider_z[63:32];
        double_divider_z_ack <= 0;
        state <= execute;
      end
    end

     double_to_long_write_a:
     begin
       double_to_long_in_stb <= 1;
       if (double_to_long_in_stb && double_to_long_in_ack) begin
         double_to_long_in_stb <= 0;
         state <= double_to_long_read_z;
       end
     end

     double_to_long_read_z:
     begin
       double_to_long_out_ack <= 1;
       if (double_to_long_out_stb && double_to_long_out_ack) begin
         double_to_long_out_ack <= 0;
         a_lo <= double_to_long_out[31:0];
         a_hi <= double_to_long_out[63:32];
         state <= execute;
       end
     end

     long_to_double_write_a:
     begin
       long_to_double_in_stb <= 1;
       if (long_to_double_in_stb && long_to_double_in_ack) begin
         long_to_double_in_stb <= 0;
         state <= long_to_double_read_z;
       end
     end

     long_to_double_read_z:
     begin
       long_to_double_out_ack <= 1;
       if (long_to_double_out_stb && long_to_double_out_ack) begin
         long_to_double_out_ack <= 0;
         a_lo <= long_to_double_out[31:0];
         a_hi <= long_to_double_out[63:32];
         state <= execute;
       end
     end

    endcase

    if (rst == 1'b1) begin
      timer <= 0;
      timer_clock <= 0;
      program_counter <= 0;
      address_z_3 <= 0;
      result <= 0;
      a = 0;
      b = 0;
      z = 0;
      state <= instruction_fetch;
      s_input_eth_in_ack <= 0;
      s_input_audio_in_ack <= 0;
      s_input_rs232_rx_ack <= 0;
      s_output_eth_out_stb <= 0;
      s_output_audio_out_stb <= 0;
      s_output_frequency_out_stb <= 0;
      s_output_samples_out_stb <= 0;
      s_output_rs232_tx_stb <= 0;
      double_divider_a_stb <= 0;
      double_divider_b_stb <= 0;
      double_divider_z_ack <= 0;
      double_to_long_in_stb <= 0;
      double_to_long_out_ack <= 0;
      long_to_double_in_stb <= 0;
      long_to_double_out_ack <= 0;
    end
  end
  assign input_eth_in_ack = s_input_eth_in_ack;
  assign input_audio_in_ack = s_input_audio_in_ack;
  assign input_rs232_rx_ack = s_input_rs232_rx_ack;
  assign output_eth_out_stb = s_output_eth_out_stb;
  assign output_eth_out = s_output_eth_out;
  assign output_audio_out_stb = s_output_audio_out_stb;
  assign output_audio_out = s_output_audio_out;
  assign output_frequency_out_stb = s_output_frequency_out_stb;
  assign output_frequency_out = s_output_frequency_out;
  assign output_samples_out_stb = s_output_samples_out_stb;
  assign output_samples_out = s_output_samples_out;
  assign output_rs232_tx_stb = s_output_rs232_tx_stb;
  assign output_rs232_tx = s_output_rs232_tx;

endmodule
