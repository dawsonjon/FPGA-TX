//name : main_0
//input : input_eth_in:16
//input : input_audio_in:16
//input : input_rs232_rx:16
//output : output_eth_out:16
//output : output_audio_out:16
//output : output_frequency_out:16
//output : output_samples_out:16
//output : output_rs232_tx:16
//source_file : /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c

///+============================================================================+
///|                                                                            |
///|                     This file was generated by Chips                       |
///|                                                                            |
///|                                  Chips                                     |
///|                                                                            |
///|                      http://github.com/dawsonjon/Chips-2.0                 |
///|                                                                            |
///|                                                             Python powered |
///+============================================================================+
module main_0(input_eth_in,input_audio_in,input_rs232_rx,input_eth_in_stb,input_audio_in_stb,input_rs232_rx_stb,output_eth_out_ack,output_audio_out_ack,output_frequency_out_ack,output_samples_out_ack,output_rs232_tx_ack,clk,rst,output_eth_out,output_audio_out,output_frequency_out,output_samples_out,output_rs232_tx,output_eth_out_stb,output_audio_out_stb,output_frequency_out_stb,output_samples_out_stb,output_rs232_tx_stb,input_eth_in_ack,input_audio_in_ack,input_rs232_rx_ack,exception);
  integer file_count;
  reg [63:0] double_divider_a;
  reg [63:0] double_divider_b;
  wire [63:0] double_divider_z;
  reg double_divider_a_stb;
  wire double_divider_a_ack;
  reg double_divider_b_stb;
  wire double_divider_b_ack;
  wire double_divider_z_stb;
  reg double_divider_z_ack;
  reg [63:0] double_to_long_in;
  wire [63:0] double_to_long_out;
  wire double_to_long_out_stb;
  reg double_to_long_out_ack;
  reg double_to_long_in_stb;
  wire double_to_long_in_ack;
  reg [63:0] long_to_double_in;
  wire [63:0] long_to_double_out;
  wire long_to_double_out_stb;
  reg long_to_double_out_ack;
  reg long_to_double_in_stb;
  wire long_to_double_in_ack;
  parameter  stop = 4'd0,
  instruction_fetch = 4'd1,
  operand_fetch = 4'd2,
  execute = 4'd3,
  load = 4'd4,
  wait_state = 4'd5,
  read = 4'd6,
  write = 4'd7,
  multiply = 4'd8,
  double_divider_write_a = 4'd9,
  double_divider_write_b = 4'd10,
  double_divider_read_z = 4'd11,
  double_to_long_write_a = 4'd12,
  double_to_long_read_z = 4'd13,
  long_to_double_write_a = 4'd14,
  long_to_double_read_z = 4'd15;
  input [31:0] input_eth_in;
  input [31:0] input_audio_in;
  input [31:0] input_rs232_rx;
  input input_eth_in_stb;
  input input_audio_in_stb;
  input input_rs232_rx_stb;
  input output_eth_out_ack;
  input output_audio_out_ack;
  input output_frequency_out_ack;
  input output_samples_out_ack;
  input output_rs232_tx_ack;
  input clk;
  input rst;
  output [31:0] output_eth_out;
  output [31:0] output_audio_out;
  output [31:0] output_frequency_out;
  output [31:0] output_samples_out;
  output [31:0] output_rs232_tx;
  output output_eth_out_stb;
  output output_audio_out_stb;
  output output_frequency_out_stb;
  output output_samples_out_stb;
  output output_rs232_tx_stb;
  output input_eth_in_ack;
  output input_audio_in_ack;
  output input_rs232_rx_ack;
  reg [31:0] timer;
  reg [63:0] timer_clock;
  reg [15:0] program_counter;
  reg [15:0] program_counter_1;
  reg [15:0] program_counter_2;
  reg [44:0] instruction;
  reg [4:0] opcode_2;
  reg [3:0] a;
  reg [3:0] b;
  reg [3:0] z;
  reg write_enable;
  reg [3:0] address_a_2;
  reg [3:0] address_b_2;
  reg [3:0] address_z_2;
  reg [3:0] address_z_3;
  reg [31:0] load_data;
  reg [31:0] write_output;
  reg [31:0] write_value;
  reg [31:0] read_input;
  reg [15:0] literal_2;
  reg [31:0] a_hi;
  reg [31:0] b_hi;
  reg [31:0] a_lo;
  reg [31:0] b_lo;
  reg [63:0] long_result;
  reg [31:0] result;
  reg [15:0] address;
  reg [31:0] data_out;
  reg [31:0] data_in;
  reg [31:0] carry;
  reg [31:0] s_output_eth_out_stb;
  reg [31:0] s_output_audio_out_stb;
  reg [31:0] s_output_frequency_out_stb;
  reg [31:0] s_output_samples_out_stb;
  reg [31:0] s_output_rs232_tx_stb;
  reg [31:0] s_output_eth_out;
  reg [31:0] s_output_audio_out;
  reg [31:0] s_output_frequency_out;
  reg [31:0] s_output_samples_out;
  reg [31:0] s_output_rs232_tx;
  reg [31:0] s_input_eth_in_ack;
  reg [31:0] s_input_audio_in_ack;
  reg [31:0] s_input_rs232_rx_ack;
  reg [15:0] state;
  output reg exception;
  reg [28:0] instructions [851:0];
  reg [31:0] memory [4096:0];
  reg [31:0] registers [15:0];
  wire [31:0] operand_a;
  wire [31:0] operand_b;
  wire [31:0] register_a;
  wire [31:0] register_b;
  wire [15:0] literal;
  wire [4:0] opcode;
  wire [3:0] address_a;
  wire [3:0] address_b;
  wire [3:0] address_z;
  wire [15:0] load_address;
  wire [15:0] store_address;
  wire [31:0] store_data;
  wire  store_enable;
  reg [31:0] product_a;
  reg [31:0] product_b;
  reg [31:0] product_c;
  reg [31:0] product_d;

  //////////////////////////////////////////////////////////////////////////////
  // Floating Point Arithmetic                                                  
  //                                                                            
  // Generate IEEE 754 single precision divider, adder and multiplier           
  //                                                                            
  double_divider double_divider_inst(
    .clk(clk),
    .rst(rst),
    .input_a(double_divider_a),
    .input_a_stb(double_divider_a_stb),
    .input_a_ack(double_divider_a_ack),
    .input_b(double_divider_b),
    .input_b_stb(double_divider_b_stb),
    .input_b_ack(double_divider_b_ack),
    .output_z(double_divider_z),
    .output_z_stb(double_divider_z_stb),
    .output_z_ack(double_divider_z_ack)
  );
  double_to_long double_to_long_inst(
    .clk(clk),
    .rst(rst),
    .input_a(double_to_long_in),
    .input_a_stb(double_to_long_in_stb),
    .input_a_ack(double_to_long_in_ack),
    .output_z(double_to_long_out),
    .output_z_stb(double_to_long_out_stb),
    .output_z_ack(double_to_long_out_ack)
  );
  long_to_double long_to_double_inst(
    .clk(clk),
    .rst(rst),
    .input_a(long_to_double_in),
    .input_a_stb(long_to_double_in_stb),
    .input_a_ack(long_to_double_in_ack),
    .output_z(long_to_double_out),
    .output_z_stb(long_to_double_out_stb),
    .output_z_ack(long_to_double_out_ack)
  );

  //////////////////////////////////////////////////////////////////////////////
  // INSTRUCTION INITIALIZATION                                                 
  //                                                                            
  // Initialise the contents of the instruction memory                          
  //
  // Intruction Set
  // ==============
  // 0 {'literal': True, 'op': 'literal'}
  // 1 {'literal': True, 'op': 'addl'}
  // 2 {'literal': False, 'op': 'store'}
  // 3 {'literal': True, 'op': 'call'}
  // 4 {'literal': False, 'op': 'stop'}
  // 5 {'literal': True, 'op': 'literal_hi'}
  // 6 {'literal': False, 'op': 'load'}
  // 7 {'literal': False, 'op': 'write'}
  // 8 {'literal': False, 'op': 'a_hi'}
  // 9 {'literal': False, 'op': 'a_lo'}
  // 10 {'literal': False, 'op': 'long_to_double'}
  // 11 {'literal': False, 'op': 'b_hi'}
  // 12 {'literal': False, 'op': 'b_lo'}
  // 13 {'literal': False, 'op': 'long_float_divide'}
  // 14 {'literal': False, 'op': 'double_to_long'}
  // 15 {'literal': False, 'op': 'read'}
  // 16 {'literal': False, 'op': 'shift_right'}
  // 17 {'literal': False, 'op': 'subtract'}
  // 18 {'literal': False, 'op': 'add'}
  // 19 {'literal': False, 'op': 'greater'}
  // 20 {'literal': True, 'op': 'jmp_if_false'}
  // 21 {'literal': True, 'op': 'goto'}
  // 22 {'literal': False, 'op': 'return'}
  // 23 {'literal': False, 'op': 'equal'}
  // 24 {'literal': False, 'op': 'multiply'}
  // 25 {'literal': False, 'op': 'greater_equal'}
  // Intructions
  // ===========
  
  initial
  begin
    instructions[0] = {5'd0, 4'd3, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 83 {'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 83, 'op': 'literal'}
    instructions[1] = {5'd0, 4'd4, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 83 {'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 83, 'op': 'literal'}
    instructions[2] = {5'd1, 4'd3, 4'd3, 16'd75};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 83 {'a': 3, 'literal': 75, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 83, 'op': 'addl'}
    instructions[3] = {5'd0, 4'd8, 4'd0, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 7 {'literal': 4, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 7, 'op': 'literal'}
    instructions[4] = {5'd0, 4'd2, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 7 {'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 7, 'op': 'literal'}
    instructions[5] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 7 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 7, 'op': 'store'}
    instructions[6] = {5'd0, 4'd8, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 9 {'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 9, 'op': 'literal'}
    instructions[7] = {5'd0, 4'd2, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 9 {'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 9, 'op': 'literal'}
    instructions[8] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 9 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 9, 'op': 'store'}
    instructions[9] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 5 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 5, 'op': 'literal'}
    instructions[10] = {5'd0, 4'd2, 4'd0, 16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 5 {'literal': 2, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 5, 'op': 'literal'}
    instructions[11] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 5 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 5, 'op': 'store'}
    instructions[12] = {5'd0, 4'd8, 4'd0, 16'd5};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 8 {'literal': 5, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 8, 'op': 'literal'}
    instructions[13] = {5'd0, 4'd2, 4'd0, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 8 {'literal': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 8, 'op': 'literal'}
    instructions[14] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 8 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 8, 'op': 'store'}
    instructions[15] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 3 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 3, 'op': 'literal'}
    instructions[16] = {5'd0, 4'd2, 4'd0, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 3 {'literal': 4, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 3, 'op': 'literal'}
    instructions[17] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 3 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 3, 'op': 'store'}
    instructions[18] = {5'd0, 4'd8, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 4 {'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 4, 'op': 'literal'}
    instructions[19] = {5'd0, 4'd2, 4'd0, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 4 {'literal': 7, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 4, 'op': 'literal'}
    instructions[20] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 4 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 4, 'op': 'store'}
    instructions[21] = {5'd0, 4'd8, 4'd0, 16'd112};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'literal': 112, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'literal'}
    instructions[22] = {5'd0, 4'd2, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'literal': 8, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'literal'}
    instructions[23] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'store'}
    instructions[24] = {5'd0, 4'd8, 4'd0, 16'd108};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'literal': 108, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'literal'}
    instructions[25] = {5'd0, 4'd2, 4'd0, 16'd9};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'literal': 9, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'literal'}
    instructions[26] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'store'}
    instructions[27] = {5'd0, 4'd8, 4'd0, 16'd97};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'literal': 97, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'literal'}
    instructions[28] = {5'd0, 4'd2, 4'd0, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'literal': 10, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'literal'}
    instructions[29] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'store'}
    instructions[30] = {5'd0, 4'd8, 4'd0, 16'd121};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'literal': 121, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'literal'}
    instructions[31] = {5'd0, 4'd2, 4'd0, 16'd11};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'literal': 11, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'literal'}
    instructions[32] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'store'}
    instructions[33] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'literal'}
    instructions[34] = {5'd0, 4'd2, 4'd0, 16'd12};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'literal': 12, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'literal'}
    instructions[35] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'store'}
    instructions[36] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'literal'}
    instructions[37] = {5'd0, 4'd2, 4'd0, 16'd13};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'literal': 13, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'literal'}
    instructions[38] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'store'}
    instructions[39] = {5'd0, 4'd8, 4'd0, 16'd103};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'literal': 103, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'literal'}
    instructions[40] = {5'd0, 4'd2, 4'd0, 16'd14};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'literal': 14, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'literal'}
    instructions[41] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'store'}
    instructions[42] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'literal'}
    instructions[43] = {5'd0, 4'd2, 4'd0, 16'd15};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'literal': 15, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'literal'}
    instructions[44] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'store'}
    instructions[45] = {5'd0, 4'd8, 4'd0, 16'd97};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'literal': 97, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'literal'}
    instructions[46] = {5'd0, 4'd2, 4'd0, 16'd16};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'literal': 16, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'literal'}
    instructions[47] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'store'}
    instructions[48] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'literal'}
    instructions[49] = {5'd0, 4'd2, 4'd0, 16'd17};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'literal': 17, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'literal'}
    instructions[50] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'store'}
    instructions[51] = {5'd0, 4'd8, 4'd0, 16'd100};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'literal': 100, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'literal'}
    instructions[52] = {5'd0, 4'd2, 4'd0, 16'd18};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'literal': 18, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'literal'}
    instructions[53] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'store'}
    instructions[54] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'literal'}
    instructions[55] = {5'd0, 4'd2, 4'd0, 16'd19};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'literal': 19, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'literal'}
    instructions[56] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'store'}
    instructions[57] = {5'd0, 4'd8, 4'd0, 16'd111};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'literal': 111, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'literal'}
    instructions[58] = {5'd0, 4'd2, 4'd0, 16'd20};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'literal': 20, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'literal'}
    instructions[59] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'store'}
    instructions[60] = {5'd0, 4'd8, 4'd0, 16'd58};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'literal': 58, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'literal'}
    instructions[61] = {5'd0, 4'd2, 4'd0, 16'd21};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'literal': 21, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'literal'}
    instructions[62] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'store'}
    instructions[63] = {5'd0, 4'd8, 4'd0, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'literal': 10, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'literal'}
    instructions[64] = {5'd0, 4'd2, 4'd0, 16'd22};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'literal': 22, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'literal'}
    instructions[65] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'store'}
    instructions[66] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'literal'}
    instructions[67] = {5'd0, 4'd2, 4'd0, 16'd23};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'literal': 23, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'literal'}
    instructions[68] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'store'}
    instructions[69] = {5'd0, 4'd8, 4'd0, 16'd99};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 99, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[70] = {5'd0, 4'd2, 4'd0, 16'd25};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 25, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[71] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'store'}
    instructions[72] = {5'd0, 4'd8, 4'd0, 16'd97};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 97, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[73] = {5'd0, 4'd2, 4'd0, 16'd26};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 26, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[74] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'store'}
    instructions[75] = {5'd0, 4'd8, 4'd0, 16'd108};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 108, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[76] = {5'd0, 4'd2, 4'd0, 16'd27};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 27, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[77] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'store'}
    instructions[78] = {5'd0, 4'd8, 4'd0, 16'd99};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 99, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[79] = {5'd0, 4'd2, 4'd0, 16'd28};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 28, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[80] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'store'}
    instructions[81] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[82] = {5'd0, 4'd2, 4'd0, 16'd29};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 29, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[83] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'store'}
    instructions[84] = {5'd0, 4'd8, 4'd0, 16'd108};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 108, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[85] = {5'd0, 4'd2, 4'd0, 16'd30};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 30, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[86] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'store'}
    instructions[87] = {5'd0, 4'd8, 4'd0, 16'd97};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 97, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[88] = {5'd0, 4'd2, 4'd0, 16'd31};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 31, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[89] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'store'}
    instructions[90] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[91] = {5'd0, 4'd2, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 32, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[92] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'store'}
    instructions[93] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[94] = {5'd0, 4'd2, 4'd0, 16'd33};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 33, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[95] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'store'}
    instructions[96] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[97] = {5'd0, 4'd2, 4'd0, 16'd34};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 34, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[98] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'store'}
    instructions[99] = {5'd0, 4'd8, 4'd0, 16'd103};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 103, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[100] = {5'd0, 4'd2, 4'd0, 16'd35};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 35, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[101] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'store'}
    instructions[102] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[103] = {5'd0, 4'd2, 4'd0, 16'd36};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 36, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[104] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'store'}
    instructions[105] = {5'd0, 4'd8, 4'd0, 16'd102};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 102, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[106] = {5'd0, 4'd2, 4'd0, 16'd37};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 37, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[107] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'store'}
    instructions[108] = {5'd0, 4'd8, 4'd0, 16'd114};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 114, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[109] = {5'd0, 4'd2, 4'd0, 16'd38};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 38, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[110] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'store'}
    instructions[111] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[112] = {5'd0, 4'd2, 4'd0, 16'd39};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 39, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[113] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'store'}
    instructions[114] = {5'd0, 4'd8, 4'd0, 16'd113};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 113, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[115] = {5'd0, 4'd2, 4'd0, 16'd40};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 40, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[116] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'store'}
    instructions[117] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[118] = {5'd0, 4'd2, 4'd0, 16'd41};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 41, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[119] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'store'}
    instructions[120] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[121] = {5'd0, 4'd2, 4'd0, 16'd42};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 42, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[122] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'store'}
    instructions[123] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[124] = {5'd0, 4'd2, 4'd0, 16'd43};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 43, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[125] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'store'}
    instructions[126] = {5'd0, 4'd8, 4'd0, 16'd99};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 99, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[127] = {5'd0, 4'd2, 4'd0, 16'd44};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 44, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[128] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'store'}
    instructions[129] = {5'd0, 4'd8, 4'd0, 16'd121};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 121, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[130] = {5'd0, 4'd2, 4'd0, 16'd45};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 45, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[131] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'store'}
    instructions[132] = {5'd0, 4'd8, 4'd0, 16'd58};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 58, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[133] = {5'd0, 4'd2, 4'd0, 16'd46};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 46, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[134] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'store'}
    instructions[135] = {5'd0, 4'd8, 4'd0, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 10, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[136] = {5'd0, 4'd2, 4'd0, 16'd47};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 47, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[137] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'store'}
    instructions[138] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[139] = {5'd0, 4'd2, 4'd0, 16'd48};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 48, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[140] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'store'}
    instructions[141] = {5'd0, 4'd8, 4'd0, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 10 {'literal': 7, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 10, 'op': 'literal'}
    instructions[142] = {5'd0, 4'd2, 4'd0, 16'd49};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 10 {'literal': 49, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 10, 'op': 'literal'}
    instructions[143] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 10 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 10, 'op': 'store'}
    instructions[144] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 4 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 4, 'op': 'literal'}
    instructions[145] = {5'd0, 4'd2, 4'd0, 16'd50};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 4 {'literal': 50, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 4, 'op': 'literal'}
    instructions[146] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 4 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 4, 'op': 'store'}
    instructions[147] = {5'd0, 4'd8, 4'd0, 16'd69};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 69, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[148] = {5'd0, 4'd2, 4'd0, 16'd51};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 51, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[149] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'store'}
    instructions[150] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[151] = {5'd0, 4'd2, 4'd0, 16'd52};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 52, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[152] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'store'}
    instructions[153] = {5'd0, 4'd8, 4'd0, 16'd116};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 116, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[154] = {5'd0, 4'd2, 4'd0, 16'd53};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 53, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[155] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'store'}
    instructions[156] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[157] = {5'd0, 4'd2, 4'd0, 16'd54};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 54, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[158] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'store'}
    instructions[159] = {5'd0, 4'd8, 4'd0, 16'd114};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 114, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[160] = {5'd0, 4'd2, 4'd0, 16'd55};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 55, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[161] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'store'}
    instructions[162] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[163] = {5'd0, 4'd2, 4'd0, 16'd56};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 56, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[164] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'store'}
    instructions[165] = {5'd0, 4'd8, 4'd0, 16'd102};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 102, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[166] = {5'd0, 4'd2, 4'd0, 16'd57};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 57, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[167] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'store'}
    instructions[168] = {5'd0, 4'd8, 4'd0, 16'd114};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 114, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[169] = {5'd0, 4'd2, 4'd0, 16'd58};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 58, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[170] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'store'}
    instructions[171] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[172] = {5'd0, 4'd2, 4'd0, 16'd59};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 59, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[173] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'store'}
    instructions[174] = {5'd0, 4'd8, 4'd0, 16'd113};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 113, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[175] = {5'd0, 4'd2, 4'd0, 16'd60};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 60, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[176] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'store'}
    instructions[177] = {5'd0, 4'd8, 4'd0, 16'd117};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 117, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[178] = {5'd0, 4'd2, 4'd0, 16'd61};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 61, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[179] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'store'}
    instructions[180] = {5'd0, 4'd8, 4'd0, 16'd101};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 101, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[181] = {5'd0, 4'd2, 4'd0, 16'd62};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 62, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[182] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'store'}
    instructions[183] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[184] = {5'd0, 4'd2, 4'd0, 16'd63};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 63, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[185] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'store'}
    instructions[186] = {5'd0, 4'd8, 4'd0, 16'd99};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 99, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[187] = {5'd0, 4'd2, 4'd0, 16'd64};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 64, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[188] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'store'}
    instructions[189] = {5'd0, 4'd8, 4'd0, 16'd121};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 121, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[190] = {5'd0, 4'd2, 4'd0, 16'd65};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 65, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[191] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'store'}
    instructions[192] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[193] = {5'd0, 4'd2, 4'd0, 16'd66};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 66, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[194] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'store'}
    instructions[195] = {5'd0, 4'd8, 4'd0, 16'd105};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 105, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[196] = {5'd0, 4'd2, 4'd0, 16'd67};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 67, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[197] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'store'}
    instructions[198] = {5'd0, 4'd8, 4'd0, 16'd110};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 110, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[199] = {5'd0, 4'd2, 4'd0, 16'd68};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 68, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[200] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'store'}
    instructions[201] = {5'd0, 4'd8, 4'd0, 16'd32};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 32, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[202] = {5'd0, 4'd2, 4'd0, 16'd69};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 69, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[203] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'store'}
    instructions[204] = {5'd0, 4'd8, 4'd0, 16'd104};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 104, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[205] = {5'd0, 4'd2, 4'd0, 16'd70};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 70, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[206] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'store'}
    instructions[207] = {5'd0, 4'd8, 4'd0, 16'd122};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 122, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[208] = {5'd0, 4'd2, 4'd0, 16'd71};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 71, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[209] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'store'}
    instructions[210] = {5'd0, 4'd8, 4'd0, 16'd58};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 58, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[211] = {5'd0, 4'd2, 4'd0, 16'd72};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 72, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[212] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'store'}
    instructions[213] = {5'd0, 4'd8, 4'd0, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 10, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[214] = {5'd0, 4'd2, 4'd0, 16'd73};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 73, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[215] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'store'}
    instructions[216] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[217] = {5'd0, 4'd2, 4'd0, 16'd74};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 74, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[218] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'store'}
    instructions[219] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 83 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 83, 'op': 'addl'}
    instructions[220] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 83 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 83, 'op': 'addl'}
    instructions[221] = {5'd3, 4'd6, 4'd0, 16'd223};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 83 {'z': 6, 'label': 223, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 83, 'op': 'call'}
    instructions[222] = {5'd4, 4'd0, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 83 {'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 83, 'op': 'stop'}
    instructions[223] = {5'd1, 4'd3, 4'd3, 16'd75};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 24 {'a': 3, 'literal': 75, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 24, 'op': 'addl'}
    instructions[224] = {5'd0, 4'd8, 4'd0, 16'd58032};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 26 {'literal': 58032, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 26, 'op': 'literal'}
    instructions[225] = {5'd5, 4'd8, 4'd8, 16'd13};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 26 {'a': 8, 'literal': 13, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 26, 'op': 'literal_hi'}
    instructions[226] = {5'd1, 4'd2, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 26 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 26, 'op': 'addl'}
    instructions[227] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 26 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 26, 'op': 'store'}
    instructions[228] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27, 'op': 'literal'}
    instructions[229] = {5'd1, 4'd2, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27 {'a': 4, 'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27, 'op': 'addl'}
    instructions[230] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27, 'op': 'store'}
    instructions[231] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27, 'op': 'literal'}
    instructions[232] = {5'd1, 4'd2, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27 {'a': 4, 'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27, 'op': 'addl'}
    instructions[233] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27, 'op': 'store'}
    instructions[234] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27, 'op': 'literal'}
    instructions[235] = {5'd1, 4'd2, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27 {'a': 4, 'literal': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27, 'op': 'addl'}
    instructions[236] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27, 'op': 'store'}
    instructions[237] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27, 'op': 'literal'}
    instructions[238] = {5'd1, 4'd2, 4'd4, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27 {'a': 4, 'literal': 4, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27, 'op': 'addl'}
    instructions[239] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27, 'op': 'store'}
    instructions[240] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27, 'op': 'literal'}
    instructions[241] = {5'd1, 4'd2, 4'd4, 16'd5};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27 {'a': 4, 'literal': 5, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27, 'op': 'addl'}
    instructions[242] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 27, 'op': 'store'}
    instructions[243] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28, 'op': 'literal'}
    instructions[244] = {5'd1, 4'd2, 4'd4, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28 {'a': 4, 'literal': 6, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28, 'op': 'addl'}
    instructions[245] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28, 'op': 'store'}
    instructions[246] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28, 'op': 'literal'}
    instructions[247] = {5'd1, 4'd2, 4'd4, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28 {'a': 4, 'literal': 7, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28, 'op': 'addl'}
    instructions[248] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28, 'op': 'store'}
    instructions[249] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28, 'op': 'literal'}
    instructions[250] = {5'd1, 4'd2, 4'd4, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28 {'a': 4, 'literal': 8, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28, 'op': 'addl'}
    instructions[251] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28, 'op': 'store'}
    instructions[252] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28, 'op': 'literal'}
    instructions[253] = {5'd1, 4'd2, 4'd4, 16'd9};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28 {'a': 4, 'literal': 9, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28, 'op': 'addl'}
    instructions[254] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28, 'op': 'store'}
    instructions[255] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28, 'op': 'literal'}
    instructions[256] = {5'd1, 4'd2, 4'd4, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28 {'a': 4, 'literal': 10, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28, 'op': 'addl'}
    instructions[257] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 28, 'op': 'store'}
    instructions[258] = {5'd0, 4'd8, 4'd0, 16'd49};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 30 {'literal': 49, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 30, 'op': 'literal'}
    instructions[259] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 30 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 30, 'op': 'addl'}
    instructions[260] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 30 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 30, 'op': 'load'}
    instructions[261] = {5'd0, 4'd2, 4'd0, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 30 {'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 30, 'op': 'literal'}
    instructions[262] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 30 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 30, 'op': 'store'}
    instructions[263] = {5'd0, 4'd8, 4'd0, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 31 {'literal': 7, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 31, 'op': 'literal'}
    instructions[264] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 31 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 31, 'op': 'addl'}
    instructions[265] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 31 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 31, 'op': 'load'}
    instructions[266] = {5'd0, 4'd2, 4'd0, 16'd50};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 31 {'literal': 50, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 31, 'op': 'literal'}
    instructions[267] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 31 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 31, 'op': 'store'}
    instructions[268] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 33 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 33, 'op': 'literal'}
    instructions[269] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 33 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 33, 'op': 'addl'}
    instructions[270] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 33 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 33, 'op': 'load'}
    instructions[271] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 33 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 33, 'op': 'store'}
    instructions[272] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 33 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 33, 'op': 'addl'}
    instructions[273] = {5'd0, 4'd8, 4'd0, 16'd16384};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 33 {'literal': 16384, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 33, 'op': 'literal'}
    instructions[274] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 33 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 33, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[275] = {5'd6, 4'd0, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 33 {'a': 3, 'z': 0, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 33, 'op': 'load'}
    instructions[276] = {5'd7, 4'd0, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 33 {'a': 0, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 33, 'op': 'write'}
    instructions[277] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 33 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 33, 'op': 'addl'}
    instructions[278] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'store'}
    instructions[279] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'addl'}
    instructions[280] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'store'}
    instructions[281] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'addl'}
    instructions[282] = {5'd0, 4'd8, 4'd0, 16'd51};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'literal': 51, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'literal'}
    instructions[283] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'store'}
    instructions[284] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'addl'}
    instructions[285] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'addl'}
    instructions[286] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'addl'}
    instructions[287] = {5'd3, 4'd6, 4'd0, 16'd584};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'z': 6, 'label': 584, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'call'}
    instructions[288] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'addl'}
    instructions[289] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[290] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'load'}
    instructions[291] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[292] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'load'}
    instructions[293] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 34, 'op': 'addl'}
    instructions[294] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35, 'op': 'store'}
    instructions[295] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35, 'op': 'addl'}
    instructions[296] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35, 'op': 'store'}
    instructions[297] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35, 'op': 'addl'}
    instructions[298] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35, 'op': 'addl'}
    instructions[299] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35, 'op': 'addl'}
    instructions[300] = {5'd3, 4'd6, 4'd0, 16'd675};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35 {'z': 6, 'label': 675, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35, 'op': 'call'}
    instructions[301] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35, 'op': 'addl'}
    instructions[302] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[303] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35, 'op': 'load'}
    instructions[304] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[305] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35, 'op': 'load'}
    instructions[306] = {5'd0, 4'd2, 4'd0, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35 {'literal': 6, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35, 'op': 'literal'}
    instructions[307] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35, 'op': 'load'}
    instructions[308] = {5'd1, 4'd2, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35, 'op': 'addl'}
    instructions[309] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 35, 'op': 'store'}
    instructions[310] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'store'}
    instructions[311] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'addl'}
    instructions[312] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'store'}
    instructions[313] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'addl'}
    instructions[314] = {5'd0, 4'd8, 4'd0, 16'd25};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'literal': 25, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'literal'}
    instructions[315] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'store'}
    instructions[316] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'addl'}
    instructions[317] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'addl'}
    instructions[318] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'addl'}
    instructions[319] = {5'd3, 4'd6, 4'd0, 16'd584};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'z': 6, 'label': 584, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'call'}
    instructions[320] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'addl'}
    instructions[321] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[322] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'load'}
    instructions[323] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[324] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'load'}
    instructions[325] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 36, 'op': 'addl'}
    instructions[326] = {5'd0, 4'd8, 4'd0, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37 {'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37, 'op': 'literal'}
    instructions[327] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37, 'op': 'addl'}
    instructions[328] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37, 'op': 'load'}
    instructions[329] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37, 'op': 'store'}
    instructions[330] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37, 'op': 'addl'}
    instructions[331] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37, 'op': 'literal'}
    instructions[332] = {5'd0, 4'd9, 4'd0, 16'd52581};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37 {'literal': 52581, 'z': 9, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37, 'op': 'literal'}
    instructions[333] = {5'd5, 4'd9, 4'd9, 16'd16333};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37 {'a': 9, 'literal': 16333, 'z': 9, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37, 'op': 'literal_hi'}
    instructions[334] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37, 'op': 'store'}
    instructions[335] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37, 'op': 'addl'}
    instructions[336] = {5'd2, 4'd0, 4'd3, 16'd9};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37 {'a': 3, 'comment': 'push', 'b': 9, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37, 'op': 'store'}
    instructions[337] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37, 'op': 'addl'}
    instructions[338] = {5'd1, 4'd8, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37, 'op': 'addl'}
    instructions[339] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37, 'op': 'addl'}
    instructions[340] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37, 'op': 'load'}
    instructions[341] = {5'd0, 4'd9, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37 {'literal': 0, 'z': 9, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37, 'op': 'literal'}
    instructions[342] = {5'd8, 4'd9, 4'd9, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37 {'a': 9, 'z': 9, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37, 'op': 'a_hi'}
    instructions[343] = {5'd9, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37 {'a': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37, 'op': 'a_lo'}
    instructions[344] = {5'd10, 4'd0, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37 {'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37, 'op': 'long_to_double'}
    instructions[345] = {5'd9, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37 {'a': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37, 'op': 'a_lo'}
    instructions[346] = {5'd8, 4'd9, 4'd9, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37 {'a': 9, 'z': 9, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37, 'op': 'a_hi'}
    instructions[347] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[348] = {5'd6, 4'd11, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37 {'a': 3, 'z': 11, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37, 'op': 'load'}
    instructions[349] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[350] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37, 'op': 'load'}
    instructions[351] = {5'd11, 4'd11, 4'd11, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37 {'a': 11, 'z': 11, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37, 'op': 'b_hi'}
    instructions[352] = {5'd12, 4'd10, 4'd10, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37 {'a': 10, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37, 'op': 'b_lo'}
    instructions[353] = {5'd8, 4'd9, 4'd9, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37 {'a': 9, 'z': 9, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37, 'op': 'a_hi'}
    instructions[354] = {5'd9, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37 {'a': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37, 'op': 'a_lo'}
    instructions[355] = {5'd13, 4'd0, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37 {'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37, 'op': 'long_float_divide'}
    instructions[356] = {5'd9, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37 {'a': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37, 'op': 'a_lo'}
    instructions[357] = {5'd8, 4'd9, 4'd9, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37 {'a': 9, 'z': 9, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37, 'op': 'a_hi'}
    instructions[358] = {5'd8, 4'd9, 4'd9, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37 {'a': 9, 'z': 9, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37, 'op': 'a_hi'}
    instructions[359] = {5'd9, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37 {'a': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37, 'op': 'a_lo'}
    instructions[360] = {5'd14, 4'd0, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37 {'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37, 'op': 'double_to_long'}
    instructions[361] = {5'd9, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37 {'a': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37, 'op': 'a_lo'}
    instructions[362] = {5'd8, 4'd9, 4'd9, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37 {'a': 9, 'z': 9, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37, 'op': 'a_hi'}
    instructions[363] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[364] = {5'd6, 4'd0, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37 {'a': 3, 'z': 0, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37, 'op': 'load'}
    instructions[365] = {5'd7, 4'd0, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37 {'a': 0, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37, 'op': 'write'}
    instructions[366] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 37, 'op': 'addl'}
    instructions[367] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'store'}
    instructions[368] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'addl'}
    instructions[369] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'store'}
    instructions[370] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'addl'}
    instructions[371] = {5'd0, 4'd8, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'literal': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'literal'}
    instructions[372] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'store'}
    instructions[373] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'addl'}
    instructions[374] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'addl'}
    instructions[375] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'addl'}
    instructions[376] = {5'd3, 4'd6, 4'd0, 16'd584};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'z': 6, 'label': 584, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'call'}
    instructions[377] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'addl'}
    instructions[378] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[379] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'load'}
    instructions[380] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[381] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'load'}
    instructions[382] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 38, 'op': 'addl'}
    instructions[383] = {5'd1, 4'd8, 4'd4, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'a': 4, 'literal': 7, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'addl'}
    instructions[384] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'addl'}
    instructions[385] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'load'}
    instructions[386] = {5'd1, 4'd2, 4'd4, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'a': 4, 'literal': 10, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'addl'}
    instructions[387] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 46, 'op': 'store'}
    instructions[388] = {5'd0, 4'd8, 4'd0, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 47 {'literal': 4, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 47, 'op': 'literal'}
    instructions[389] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 47 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 47, 'op': 'addl'}
    instructions[390] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 47 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 47, 'op': 'load'}
    instructions[391] = {5'd15, 4'd8, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 47 {'a': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 47, 'op': 'read'}
    instructions[392] = {5'd1, 4'd2, 4'd4, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 47 {'a': 4, 'literal': 7, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 47, 'op': 'addl'}
    instructions[393] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 47 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 47, 'op': 'store'}
    instructions[394] = {5'd0, 4'd8, 4'd0, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 48 {'literal': 10, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 48, 'op': 'literal'}
    instructions[395] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 48 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 48, 'op': 'store'}
    instructions[396] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 48 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 48, 'op': 'addl'}
    instructions[397] = {5'd1, 4'd8, 4'd4, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 48 {'a': 4, 'literal': 7, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 48, 'op': 'addl'}
    instructions[398] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 48 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 48, 'op': 'addl'}
    instructions[399] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 48 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 48, 'op': 'load'}
    instructions[400] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 48 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 48, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[401] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 48 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 48, 'op': 'load'}
    instructions[402] = {5'd16, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 48 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 48, 'op': 'shift_right'}
    instructions[403] = {5'd1, 4'd2, 4'd4, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 48 {'a': 4, 'literal': 7, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 48, 'op': 'addl'}
    instructions[404] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 48 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 48, 'op': 'store'}
    instructions[405] = {5'd1, 4'd8, 4'd4, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 49 {'a': 4, 'literal': 10, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 49, 'op': 'addl'}
    instructions[406] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 49 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 49, 'op': 'addl'}
    instructions[407] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 49 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 49, 'op': 'load'}
    instructions[408] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 49 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 49, 'op': 'store'}
    instructions[409] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 49 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 49, 'op': 'addl'}
    instructions[410] = {5'd1, 4'd8, 4'd4, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 49 {'a': 4, 'literal': 7, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 49, 'op': 'addl'}
    instructions[411] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 49 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 49, 'op': 'addl'}
    instructions[412] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 49 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 49, 'op': 'load'}
    instructions[413] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 49 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 49, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[414] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 49 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 49, 'op': 'load'}
    instructions[415] = {5'd17, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 49 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 49, 'op': 'subtract'}
    instructions[416] = {5'd1, 4'd2, 4'd4, 16'd5};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 49 {'a': 4, 'literal': 5, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 49, 'op': 'addl'}
    instructions[417] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 49 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 49, 'op': 'store'}
    instructions[418] = {5'd1, 4'd8, 4'd4, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 52 {'a': 4, 'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 52, 'op': 'addl'}
    instructions[419] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 52 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 52, 'op': 'addl'}
    instructions[420] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 52 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 52, 'op': 'load'}
    instructions[421] = {5'd1, 4'd2, 4'd4, 16'd9};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 52 {'a': 4, 'literal': 9, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 52, 'op': 'addl'}
    instructions[422] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 52 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 52, 'op': 'store'}
    instructions[423] = {5'd1, 4'd8, 4'd4, 16'd5};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 54 {'a': 4, 'literal': 5, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 54, 'op': 'addl'}
    instructions[424] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 54 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 54, 'op': 'addl'}
    instructions[425] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 54 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 54, 'op': 'load'}
    instructions[426] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 54 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 54, 'op': 'store'}
    instructions[427] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 54 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 54, 'op': 'addl'}
    instructions[428] = {5'd1, 4'd8, 4'd4, 16'd9};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 54 {'a': 4, 'literal': 9, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 54, 'op': 'addl'}
    instructions[429] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 54 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 54, 'op': 'addl'}
    instructions[430] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 54 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 54, 'op': 'load'}
    instructions[431] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 54 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 54, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[432] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 54 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 54, 'op': 'load'}
    instructions[433] = {5'd18, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 54 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 54, 'op': 'add'}
    instructions[434] = {5'd1, 4'd2, 4'd4, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 54 {'a': 4, 'literal': 6, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 54, 'op': 'addl'}
    instructions[435] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 54 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 54, 'op': 'store'}
    instructions[436] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57, 'op': 'addl'}
    instructions[437] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57, 'op': 'addl'}
    instructions[438] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57, 'op': 'load'}
    instructions[439] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57, 'op': 'store'}
    instructions[440] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57, 'op': 'addl'}
    instructions[441] = {5'd1, 4'd8, 4'd4, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57 {'a': 4, 'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57, 'op': 'addl'}
    instructions[442] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57, 'op': 'addl'}
    instructions[443] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57, 'op': 'load'}
    instructions[444] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[445] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57, 'op': 'load'}
    instructions[446] = {5'd19, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57, 'op': 'greater'}
    instructions[447] = {5'd20, 4'd0, 4'd8, 16'd454};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57 {'a': 8, 'label': 454, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57, 'op': 'jmp_if_false'}
    instructions[448] = {5'd1, 4'd8, 4'd4, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57 {'a': 4, 'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57, 'op': 'addl'}
    instructions[449] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57, 'op': 'addl'}
    instructions[450] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57, 'op': 'load'}
    instructions[451] = {5'd1, 4'd2, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57 {'a': 4, 'literal': 2, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57, 'op': 'addl'}
    instructions[452] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57, 'op': 'store'}
    instructions[453] = {5'd21, 4'd0, 4'd0, 16'd454};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57 {'label': 454, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 57, 'op': 'goto'}
    instructions[454] = {5'd1, 4'd8, 4'd4, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 58 {'a': 4, 'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 58, 'op': 'addl'}
    instructions[455] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 58 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 58, 'op': 'addl'}
    instructions[456] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 58 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 58, 'op': 'load'}
    instructions[457] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 58 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 58, 'op': 'store'}
    instructions[458] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 58 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 58, 'op': 'addl'}
    instructions[459] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 58 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 58, 'op': 'addl'}
    instructions[460] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 58 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 58, 'op': 'addl'}
    instructions[461] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 58 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 58, 'op': 'load'}
    instructions[462] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 58 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 58, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[463] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 58 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 58, 'op': 'load'}
    instructions[464] = {5'd19, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 58 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 58, 'op': 'greater'}
    instructions[465] = {5'd20, 4'd0, 4'd8, 16'd472};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 58 {'a': 8, 'label': 472, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 58, 'op': 'jmp_if_false'}
    instructions[466] = {5'd1, 4'd8, 4'd4, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 58 {'a': 4, 'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 58, 'op': 'addl'}
    instructions[467] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 58 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 58, 'op': 'addl'}
    instructions[468] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 58 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 58, 'op': 'load'}
    instructions[469] = {5'd1, 4'd2, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 58 {'a': 4, 'literal': 1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 58, 'op': 'addl'}
    instructions[470] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 58 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 58, 'op': 'store'}
    instructions[471] = {5'd21, 4'd0, 4'd0, 16'd472};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 58 {'label': 472, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 58, 'op': 'goto'}
    instructions[472] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 59 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 59, 'op': 'literal'}
    instructions[473] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 59 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 59, 'op': 'store'}
    instructions[474] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 59 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 59, 'op': 'addl'}
    instructions[475] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 59 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 59, 'op': 'addl'}
    instructions[476] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 59 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 59, 'op': 'addl'}
    instructions[477] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 59 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 59, 'op': 'load'}
    instructions[478] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 59 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 59, 'op': 'store'}
    instructions[479] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 59 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 59, 'op': 'addl'}
    instructions[480] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 59 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 59, 'op': 'addl'}
    instructions[481] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 59 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 59, 'op': 'addl'}
    instructions[482] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 59 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 59, 'op': 'load'}
    instructions[483] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 59 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 59, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[484] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 59 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 59, 'op': 'load'}
    instructions[485] = {5'd18, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 59 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 59, 'op': 'add'}
    instructions[486] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 59 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 59, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[487] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 59 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 59, 'op': 'load'}
    instructions[488] = {5'd16, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 59 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 59, 'op': 'shift_right'}
    instructions[489] = {5'd1, 4'd2, 4'd4, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 59 {'a': 4, 'literal': 8, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 59, 'op': 'addl'}
    instructions[490] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 59 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 59, 'op': 'store'}
    instructions[491] = {5'd1, 4'd8, 4'd4, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 60 {'a': 4, 'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 60, 'op': 'addl'}
    instructions[492] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 60 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 60, 'op': 'addl'}
    instructions[493] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 60 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 60, 'op': 'load'}
    instructions[494] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 60 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 60, 'op': 'store'}
    instructions[495] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 60 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 60, 'op': 'addl'}
    instructions[496] = {5'd1, 4'd8, 4'd4, 16'd2};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 60 {'a': 4, 'literal': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 60, 'op': 'addl'}
    instructions[497] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 60 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 60, 'op': 'addl'}
    instructions[498] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 60 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 60, 'op': 'load'}
    instructions[499] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 60 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 60, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[500] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 60 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 60, 'op': 'load'}
    instructions[501] = {5'd17, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 60 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 60, 'op': 'subtract'}
    instructions[502] = {5'd1, 4'd2, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 60 {'a': 4, 'literal': 3, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 60, 'op': 'addl'}
    instructions[503] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 60 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 60, 'op': 'store'}
    instructions[504] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 61 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 61, 'op': 'literal'}
    instructions[505] = {5'd1, 4'd2, 4'd4, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 61 {'a': 4, 'literal': 4, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 61, 'op': 'addl'}
    instructions[506] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 61 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 61, 'op': 'store'}
    instructions[507] = {5'd0, 4'd8, 4'd0, 16'd256};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 62 {'literal': 256, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 62, 'op': 'literal'}
    instructions[508] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 62 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 62, 'op': 'store'}
    instructions[509] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 62 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 62, 'op': 'addl'}
    instructions[510] = {5'd1, 4'd8, 4'd4, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 62 {'a': 4, 'literal': 4, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 62, 'op': 'addl'}
    instructions[511] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 62 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 62, 'op': 'addl'}
    instructions[512] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 62 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 62, 'op': 'load'}
    instructions[513] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 62 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 62, 'op': 'store'}
    instructions[514] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 62 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 62, 'op': 'addl'}
    instructions[515] = {5'd1, 4'd8, 4'd4, 16'd3};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 62 {'a': 4, 'literal': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 62, 'op': 'addl'}
    instructions[516] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 62 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 62, 'op': 'addl'}
    instructions[517] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 62 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 62, 'op': 'load'}
    instructions[518] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 62 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 62, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[519] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 62 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 62, 'op': 'load'}
    instructions[520] = {5'd16, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 62 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 62, 'op': 'shift_right'}
    instructions[521] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 62 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 62, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[522] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 62 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 62, 'op': 'load'}
    instructions[523] = {5'd19, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 62 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 62, 'op': 'greater'}
    instructions[524] = {5'd20, 4'd0, 4'd8, 16'd544};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 8, 'label': 544, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'jmp_if_false'}
    instructions[525] = {5'd1, 4'd8, 4'd4, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 63 {'a': 4, 'literal': 4, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 63, 'op': 'addl'}
    instructions[526] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 63 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 63, 'op': 'addl'}
    instructions[527] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 63 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 63, 'op': 'load'}
    instructions[528] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 63 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 63, 'op': 'store'}
    instructions[529] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 63 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 63, 'op': 'addl'}
    instructions[530] = {5'd0, 4'd8, 4'd0, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 63 {'literal': 1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 63, 'op': 'literal'}
    instructions[531] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 63 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 63, 'op': 'store'}
    instructions[532] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 63 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 63, 'op': 'addl'}
    instructions[533] = {5'd1, 4'd8, 4'd4, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 63 {'a': 4, 'literal': 4, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 63, 'op': 'addl'}
    instructions[534] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 63 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 63, 'op': 'addl'}
    instructions[535] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 63 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 63, 'op': 'load'}
    instructions[536] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 63 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 63, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[537] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 63 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 63, 'op': 'load'}
    instructions[538] = {5'd18, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 63 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 63, 'op': 'add'}
    instructions[539] = {5'd1, 4'd2, 4'd4, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 63 {'a': 4, 'literal': 4, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 63, 'op': 'addl'}
    instructions[540] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 63 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 63, 'op': 'store'}
    instructions[541] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 63 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 63, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[542] = {5'd6, 4'd8, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 63 {'a': 3, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 63, 'op': 'load'}
    instructions[543] = {5'd21, 4'd0, 4'd0, 16'd545};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'label': 545, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'goto'}
    instructions[544] = {5'd21, 4'd0, 4'd0, 16'd546};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'label': 546, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'goto'}
    instructions[545] = {5'd21, 4'd0, 4'd0, 16'd507};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 62 {'label': 507, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 62, 'op': 'goto'}
    instructions[546] = {5'd2, 4'd0, 4'd3, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'store'}
    instructions[547] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'addl'}
    instructions[548] = {5'd2, 4'd0, 4'd3, 16'd7};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'store'}
    instructions[549] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'addl'}
    instructions[550] = {5'd1, 4'd8, 4'd4, 16'd4};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 4, 'literal': 4, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'addl'}
    instructions[551] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'addl'}
    instructions[552] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'load'}
    instructions[553] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'store'}
    instructions[554] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'addl'}
    instructions[555] = {5'd1, 4'd8, 4'd4, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 4, 'literal': 8, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'addl'}
    instructions[556] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'addl'}
    instructions[557] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'load'}
    instructions[558] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'store'}
    instructions[559] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'addl'}
    instructions[560] = {5'd1, 4'd8, 4'd4, 16'd6};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 4, 'literal': 6, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'addl'}
    instructions[561] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'addl'}
    instructions[562] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'load'}
    instructions[563] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[564] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'load'}
    instructions[565] = {5'd17, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'subtract'}
    instructions[566] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[567] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'load'}
    instructions[568] = {5'd16, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'shift_right'}
    instructions[569] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'store'}
    instructions[570] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'addl'}
    instructions[571] = {5'd1, 4'd7, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'addl'}
    instructions[572] = {5'd1, 4'd4, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'addl'}
    instructions[573] = {5'd3, 4'd6, 4'd0, 16'd802};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'z': 6, 'label': 802, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'call'}
    instructions[574] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 3, 'literal': -1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'addl'}
    instructions[575] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[576] = {5'd6, 4'd7, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 3, 'z': 7, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'load'}
    instructions[577] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[578] = {5'd6, 4'd6, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 3, 'z': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'load'}
    instructions[579] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 65, 'op': 'addl'}
    instructions[580] = {5'd21, 4'd0, 4'd0, 16'd383};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 40 {'label': 383, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 40, 'op': 'goto'}
    instructions[581] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 24 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 24, 'op': 'addl'}
    instructions[582] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 24 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 24, 'op': 'addl'}
    instructions[583] = {5'd22, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 24 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 24, 'op': 'return'}
    instructions[584] = {5'd1, 4'd3, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73 {'a': 3, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73, 'op': 'addl'}
    instructions[585] = {5'd2, 4'd0, 4'd3, 16'd6};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'store'}
    instructions[586] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[587] = {5'd2, 4'd0, 4'd3, 16'd7};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'store'}
    instructions[588] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[589] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[590] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[591] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'load'}
    instructions[592] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'store'}
    instructions[593] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[594] = {5'd0, 4'd8, 4'd0, 16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'literal': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'literal'}
    instructions[595] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[596] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'load'}
    instructions[597] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'store'}
    instructions[598] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[599] = {5'd1, 4'd7, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 4, 'literal': 0, 'z': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[600] = {5'd1, 4'd4, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[601] = {5'd3, 4'd6, 4'd0, 16'd611};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'z': 6, 'label': 611, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'call'}
    instructions[602] = {5'd1, 4'd3, 4'd3, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': -2, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[603] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[604] = {5'd6, 4'd7, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'z': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'load'}
    instructions[605] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[606] = {5'd6, 4'd6, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'z': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'load'}
    instructions[607] = {5'd1, 4'd3, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74 {'a': 3, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 74, 'op': 'addl'}
    instructions[608] = {5'd1, 4'd3, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73 {'a': 4, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73, 'op': 'addl'}
    instructions[609] = {5'd1, 4'd4, 4'd7, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73 {'a': 7, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73, 'op': 'addl'}
    instructions[610] = {5'd22, 4'd0, 4'd6, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73 {'a': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 73, 'op': 'return'}
    instructions[611] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23, 'op': 'addl'}
    instructions[612] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 24 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 24, 'op': 'literal'}
    instructions[613] = {5'd1, 4'd2, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 24 {'a': 4, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 24, 'op': 'addl'}
    instructions[614] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 24 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 24, 'op': 'store'}
    instructions[615] = {5'd1, 4'd8, 4'd4, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 4, 'literal': -2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'addl'}
    instructions[616] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'addl'}
    instructions[617] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'load'}
    instructions[618] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'store'}
    instructions[619] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'addl'}
    instructions[620] = {5'd1, 4'd8, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 4, 'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'addl'}
    instructions[621] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'addl'}
    instructions[622] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'load'}
    instructions[623] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[624] = {5'd6, 4'd2, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 3, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'load'}
    instructions[625] = {5'd18, 4'd8, 4'd8, 16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 8, 'z': 8, 'b': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'add'}
    instructions[626] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'addl'}
    instructions[627] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'load'}
    instructions[628] = {5'd20, 4'd0, 4'd8, 16'd670};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 29 {'a': 8, 'label': 670, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 29, 'op': 'jmp_if_false'}
    instructions[629] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[630] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[631] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'load'}
    instructions[632] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'store'}
    instructions[633] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[634] = {5'd1, 4'd8, 4'd4, -16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 4, 'literal': -2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[635] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[636] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'load'}
    instructions[637] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'store'}
    instructions[638] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[639] = {5'd1, 4'd8, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 4, 'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[640] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[641] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'load'}
    instructions[642] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[643] = {5'd6, 4'd2, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'load'}
    instructions[644] = {5'd18, 4'd8, 4'd8, 16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 8, 'z': 8, 'b': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'add'}
    instructions[645] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[646] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'load'}
    instructions[647] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[648] = {5'd6, 4'd0, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'z': 0, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'load'}
    instructions[649] = {5'd7, 4'd0, 4'd0, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 0, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'write'}
    instructions[650] = {5'd1, 4'd3, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26 {'a': 3, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 26, 'op': 'addl'}
    instructions[651] = {5'd1, 4'd8, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 4, 'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[652] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[653] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'load'}
    instructions[654] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'store'}
    instructions[655] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[656] = {5'd0, 4'd8, 4'd0, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'literal': 1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'literal'}
    instructions[657] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'store'}
    instructions[658] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[659] = {5'd1, 4'd8, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 4, 'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[660] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[661] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'load'}
    instructions[662] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[663] = {5'd6, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'load'}
    instructions[664] = {5'd18, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'add'}
    instructions[665] = {5'd1, 4'd2, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 4, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'addl'}
    instructions[666] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'store'}
    instructions[667] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[668] = {5'd6, 4'd8, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27 {'a': 3, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 27, 'op': 'load'}
    instructions[669] = {5'd21, 4'd0, 4'd0, 16'd671};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 29 {'label': 671, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 29, 'op': 'goto'}
    instructions[670] = {5'd21, 4'd0, 4'd0, 16'd672};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 29 {'label': 672, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 29, 'op': 'goto'}
    instructions[671] = {5'd21, 4'd0, 4'd0, 16'd615};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25 {'label': 615, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 25, 'op': 'goto'}
    instructions[672] = {5'd1, 4'd3, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23 {'a': 4, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23, 'op': 'addl'}
    instructions[673] = {5'd1, 4'd4, 4'd7, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23 {'a': 7, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23, 'op': 'addl'}
    instructions[674] = {5'd22, 4'd0, 4'd6, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23 {'a': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/stdio.h : 23, 'op': 'return'}
    instructions[675] = {5'd1, 4'd3, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 155 {'a': 3, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 155, 'op': 'addl'}
    instructions[676] = {5'd2, 4'd0, 4'd3, 16'd6};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'op': 'store'}
    instructions[677] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'op': 'addl'}
    instructions[678] = {5'd2, 4'd0, 4'd3, 16'd7};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'op': 'store'}
    instructions[679] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'op': 'addl'}
    instructions[680] = {5'd0, 4'd8, 4'd0, 16'd50};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'literal': 50, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'op': 'literal'}
    instructions[681] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'op': 'addl'}
    instructions[682] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'op': 'load'}
    instructions[683] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'op': 'store'}
    instructions[684] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'op': 'addl'}
    instructions[685] = {5'd1, 4'd7, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'a': 4, 'literal': 0, 'z': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'op': 'addl'}
    instructions[686] = {5'd1, 4'd4, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'a': 3, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'op': 'addl'}
    instructions[687] = {5'd3, 4'd6, 4'd0, 16'd700};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'z': 6, 'label': 700, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'op': 'call'}
    instructions[688] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'a': 3, 'literal': -1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'op': 'addl'}
    instructions[689] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[690] = {5'd6, 4'd7, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'a': 3, 'z': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'op': 'load'}
    instructions[691] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[692] = {5'd6, 4'd6, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'a': 3, 'z': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'op': 'load'}
    instructions[693] = {5'd0, 4'd2, 4'd0, 16'd5};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'literal': 5, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'op': 'literal'}
    instructions[694] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'op': 'load'}
    instructions[695] = {5'd0, 4'd2, 4'd0, 16'd6};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'literal': 6, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'op': 'literal'}
    instructions[696] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'op': 'store'}
    instructions[697] = {5'd1, 4'd3, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'a': 4, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'op': 'addl'}
    instructions[698] = {5'd1, 4'd4, 4'd7, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'a': 7, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'op': 'addl'}
    instructions[699] = {5'd22, 4'd0, 4'd6, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156 {'a': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 156, 'op': 'return'}
    instructions[700] = {5'd1, 4'd3, 4'd3, 16'd2};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 26 {'a': 3, 'literal': 2, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 26, 'op': 'addl'}
    instructions[701] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 29 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 29, 'op': 'literal'}
    instructions[702] = {5'd1, 4'd2, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 29 {'a': 4, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 29, 'op': 'addl'}
    instructions[703] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 29 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 29, 'op': 'store'}
    instructions[704] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 31 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 31, 'op': 'addl'}
    instructions[705] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 31 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 31, 'op': 'addl'}
    instructions[706] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 31 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 31, 'op': 'load'}
    instructions[707] = {5'd15, 4'd8, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 31 {'a': 8, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 31, 'op': 'read'}
    instructions[708] = {5'd1, 4'd2, 4'd4, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 31 {'a': 4, 'literal': 1, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 31, 'op': 'addl'}
    instructions[709] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 31 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 31, 'op': 'store'}
    instructions[710] = {5'd0, 4'd8, 4'd0, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'literal'}
    instructions[711] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'store'}
    instructions[712] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'addl'}
    instructions[713] = {5'd2, 4'd0, 4'd3, 16'd6};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'a': 3, 'comment': 'push', 'b': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'store'}
    instructions[714] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'addl'}
    instructions[715] = {5'd2, 4'd0, 4'd3, 16'd7};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'a': 3, 'comment': 'push', 'b': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'store'}
    instructions[716] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'addl'}
    instructions[717] = {5'd1, 4'd8, 4'd4, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'a': 4, 'literal': 1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'addl'}
    instructions[718] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'addl'}
    instructions[719] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'load'}
    instructions[720] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'store'}
    instructions[721] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'addl'}
    instructions[722] = {5'd1, 4'd7, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'a': 4, 'literal': 0, 'z': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'addl'}
    instructions[723] = {5'd1, 4'd4, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'a': 3, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'addl'}
    instructions[724] = {5'd3, 4'd6, 4'd0, 16'd777};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'z': 6, 'label': 777, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'call'}
    instructions[725] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'a': 3, 'literal': -1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'addl'}
    instructions[726] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[727] = {5'd6, 4'd7, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'a': 3, 'z': 7, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'load'}
    instructions[728] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[729] = {5'd6, 4'd6, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'a': 3, 'z': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'load'}
    instructions[730] = {5'd0, 4'd2, 4'd0, 16'd24};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'literal': 24, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'literal'}
    instructions[731] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'load'}
    instructions[732] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[733] = {5'd6, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'load'}
    instructions[734] = {5'd23, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'equal'}
    instructions[735] = {5'd20, 4'd0, 4'd8, 16'd738};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'a': 8, 'label': 738, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'jmp_if_false'}
    instructions[736] = {5'd21, 4'd0, 4'd0, 16'd769};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'label': 769, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'goto'}
    instructions[737] = {5'd21, 4'd0, 4'd0, 16'd738};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32 {'label': 738, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 32, 'op': 'goto'}
    instructions[738] = {5'd0, 4'd8, 4'd0, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 33 {'literal': 10, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 33, 'op': 'literal'}
    instructions[739] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 33 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 33, 'op': 'store'}
    instructions[740] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 33 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 33, 'op': 'addl'}
    instructions[741] = {5'd1, 4'd8, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 33 {'a': 4, 'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 33, 'op': 'addl'}
    instructions[742] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 33 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 33, 'op': 'addl'}
    instructions[743] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 33 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 33, 'op': 'load'}
    instructions[744] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 33 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 33, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[745] = {5'd6, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 33 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 33, 'op': 'load'}
    instructions[746] = {5'd24, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 33 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 33, 'op': 'multiply'}
    instructions[747] = {5'd1, 4'd2, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 33 {'a': 4, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 33, 'op': 'addl'}
    instructions[748] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 33 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 33, 'op': 'store'}
    instructions[749] = {5'd0, 4'd8, 4'd0, 16'd48};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34 {'literal': 48, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34, 'op': 'literal'}
    instructions[750] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34, 'op': 'store'}
    instructions[751] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34, 'op': 'addl'}
    instructions[752] = {5'd1, 4'd8, 4'd4, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34 {'a': 4, 'literal': 1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34, 'op': 'addl'}
    instructions[753] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34, 'op': 'addl'}
    instructions[754] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34, 'op': 'load'}
    instructions[755] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[756] = {5'd6, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34, 'op': 'load'}
    instructions[757] = {5'd17, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34, 'op': 'subtract'}
    instructions[758] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34, 'op': 'store'}
    instructions[759] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34, 'op': 'addl'}
    instructions[760] = {5'd1, 4'd8, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34 {'a': 4, 'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34, 'op': 'addl'}
    instructions[761] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34, 'op': 'addl'}
    instructions[762] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34, 'op': 'load'}
    instructions[763] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[764] = {5'd6, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34, 'op': 'load'}
    instructions[765] = {5'd18, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34, 'op': 'add'}
    instructions[766] = {5'd1, 4'd2, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34 {'a': 4, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34, 'op': 'addl'}
    instructions[767] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 34, 'op': 'store'}
    instructions[768] = {5'd21, 4'd0, 4'd0, 16'd704};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 30 {'label': 704, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 30, 'op': 'goto'}
    instructions[769] = {5'd1, 4'd8, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 36 {'a': 4, 'literal': 0, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 36, 'op': 'addl'}
    instructions[770] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 36 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 36, 'op': 'addl'}
    instructions[771] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 36 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 36, 'op': 'load'}
    instructions[772] = {5'd0, 4'd2, 4'd0, 16'd5};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 36 {'literal': 5, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 36, 'op': 'literal'}
    instructions[773] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 36 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 36, 'op': 'store'}
    instructions[774] = {5'd1, 4'd3, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 36 {'a': 4, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 36, 'op': 'addl'}
    instructions[775] = {5'd1, 4'd4, 4'd7, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 36 {'a': 7, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 36, 'op': 'addl'}
    instructions[776] = {5'd22, 4'd0, 4'd6, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 36 {'a': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/scan.h : 36, 'op': 'return'}
    instructions[777] = {5'd1, 4'd3, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 86 {'a': 3, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 86, 'op': 'addl'}
    instructions[778] = {5'd0, 4'd8, 4'd0, 16'd48};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'literal': 48, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'op': 'literal'}
    instructions[779] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'op': 'store'}
    instructions[780] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'op': 'addl'}
    instructions[781] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'op': 'addl'}
    instructions[782] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'op': 'addl'}
    instructions[783] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'op': 'load'}
    instructions[784] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[785] = {5'd6, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'op': 'load'}
    instructions[786] = {5'd25, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'op': 'greater_equal'}
    instructions[787] = {5'd20, 4'd0, 4'd8, 16'd797};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'a': 8, 'label': 797, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'op': 'jmp_if_false'}
    instructions[788] = {5'd1, 4'd8, 4'd4, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'a': 4, 'literal': -1, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'op': 'addl'}
    instructions[789] = {5'd1, 4'd2, 4'd8, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'a': 8, 'literal': 0, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'op': 'addl'}
    instructions[790] = {5'd6, 4'd8, 4'd2, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'a': 2, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'op': 'load'}
    instructions[791] = {5'd2, 4'd0, 4'd3, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'op': 'store'}
    instructions[792] = {5'd1, 4'd3, 4'd3, 16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'a': 3, 'literal': 1, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'op': 'addl'}
    instructions[793] = {5'd0, 4'd8, 4'd0, 16'd57};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'literal': 57, 'z': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'op': 'literal'}
    instructions[794] = {5'd1, 4'd3, 4'd3, -16'd1};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'a': 3, 'comment': 'pop', 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[795] = {5'd6, 4'd10, 4'd3, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'a': 3, 'z': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'op': 'load'}
    instructions[796] = {5'd25, 4'd8, 4'd8, 16'd10};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'a': 8, 'z': 8, 'b': 10, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'op': 'greater_equal'}
    instructions[797] = {5'd0, 4'd2, 4'd0, 16'd24};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'literal': 24, 'z': 2, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'op': 'literal'}
    instructions[798] = {5'd2, 4'd0, 4'd2, 16'd8};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'a': 2, 'b': 8, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'op': 'store'}
    instructions[799] = {5'd1, 4'd3, 4'd4, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'a': 4, 'literal': 0, 'z': 3, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'op': 'addl'}
    instructions[800] = {5'd1, 4'd4, 4'd7, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'a': 7, 'literal': 0, 'z': 4, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'op': 'addl'}
    instructions[801] = {5'd22, 4'd0, 4'd6, 16'd0};///usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87 {'a': 6, 'trace': /usr/local/lib/python2.7/dist-packages/chips/compiler/include/ctype.h : 87, 'op': 'return'}
    instructions[802] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 18 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 18, 'op': 'addl'}
    instructions[803] = {5'd0, 4'd8, 4'd0, 16'd127};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 19 {'literal': 127, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 19, 'op': 'literal'}
    instructions[804] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 19 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 19, 'op': 'store'}
    instructions[805] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 19 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 19, 'op': 'addl'}
    instructions[806] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 19 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 19, 'op': 'addl'}
    instructions[807] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 19 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 19, 'op': 'addl'}
    instructions[808] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 19 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 19, 'op': 'load'}
    instructions[809] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 19 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 19, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[810] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 19 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 19, 'op': 'load'}
    instructions[811] = {5'd19, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 19 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 19, 'op': 'greater'}
    instructions[812] = {5'd20, 4'd0, 4'd8, 16'd817};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 19 {'a': 8, 'label': 817, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 19, 'op': 'jmp_if_false'}
    instructions[813] = {5'd0, 4'd8, 4'd0, 16'd127};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 19 {'literal': 127, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 19, 'op': 'literal'}
    instructions[814] = {5'd1, 4'd2, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 19 {'a': 4, 'literal': -1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 19, 'op': 'addl'}
    instructions[815] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 19 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 19, 'op': 'store'}
    instructions[816] = {5'd21, 4'd0, 4'd0, 16'd817};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 19 {'label': 817, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 19, 'op': 'goto'}
    instructions[817] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 20 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 20, 'op': 'addl'}
    instructions[818] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 20 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 20, 'op': 'addl'}
    instructions[819] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 20 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 20, 'op': 'load'}
    instructions[820] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 20 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 20, 'op': 'store'}
    instructions[821] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 20 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 20, 'op': 'addl'}
    instructions[822] = {5'd0, 4'd8, 4'd0, 16'd65408};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 20 {'literal': 65408, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 20, 'op': 'literal'}
    instructions[823] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 20 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 20, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[824] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 20 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 20, 'op': 'load'}
    instructions[825] = {5'd19, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 20 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 20, 'op': 'greater'}
    instructions[826] = {5'd20, 4'd0, 4'd8, 16'd831};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 20 {'a': 8, 'label': 831, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 20, 'op': 'jmp_if_false'}
    instructions[827] = {5'd0, 4'd8, 4'd0, 16'd65408};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 20 {'literal': 65408, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 20, 'op': 'literal'}
    instructions[828] = {5'd1, 4'd2, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 20 {'a': 4, 'literal': -1, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 20, 'op': 'addl'}
    instructions[829] = {5'd2, 4'd0, 4'd2, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 20 {'a': 2, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 20, 'op': 'store'}
    instructions[830] = {5'd21, 4'd0, 4'd0, 16'd831};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 20 {'label': 831, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 20, 'op': 'goto'}
    instructions[831] = {5'd0, 4'd8, 4'd0, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 21 {'literal': 0, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 21, 'op': 'literal'}
    instructions[832] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 21 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 21, 'op': 'addl'}
    instructions[833] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 21 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 21, 'op': 'load'}
    instructions[834] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 21 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 21, 'op': 'store'}
    instructions[835] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 21 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 21, 'op': 'addl'}
    instructions[836] = {5'd0, 4'd8, 4'd0, 16'd128};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 21 {'literal': 128, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 21, 'op': 'literal'}
    instructions[837] = {5'd2, 4'd0, 4'd3, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 21 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 21, 'op': 'store'}
    instructions[838] = {5'd1, 4'd3, 4'd3, 16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 21 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 21, 'op': 'addl'}
    instructions[839] = {5'd1, 4'd8, 4'd4, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 21 {'a': 4, 'literal': -1, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 21, 'op': 'addl'}
    instructions[840] = {5'd1, 4'd2, 4'd8, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 21 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 21, 'op': 'addl'}
    instructions[841] = {5'd6, 4'd8, 4'd2, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 21 {'a': 2, 'z': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 21, 'op': 'load'}
    instructions[842] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 21 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 21, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[843] = {5'd6, 4'd10, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 21 {'a': 3, 'z': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 21, 'op': 'load'}
    instructions[844] = {5'd18, 4'd8, 4'd8, 16'd10};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 21 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 21, 'op': 'add'}
    instructions[845] = {5'd1, 4'd3, 4'd3, -16'd1};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 21 {'a': 3, 'comment': 'pop', 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 21, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[846] = {5'd6, 4'd0, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 21 {'a': 3, 'z': 0, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 21, 'op': 'load'}
    instructions[847] = {5'd7, 4'd0, 4'd0, 16'd8};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 21 {'a': 0, 'b': 8, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 21, 'op': 'write'}
    instructions[848] = {5'd1, 4'd3, 4'd3, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 21 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 21, 'op': 'addl'}
    instructions[849] = {5'd1, 4'd3, 4'd4, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 18 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 18, 'op': 'addl'}
    instructions[850] = {5'd1, 4'd4, 4'd7, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 18 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 18, 'op': 'addl'}
    instructions[851] = {5'd22, 4'd0, 4'd6, 16'd0};///home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 18 {'a': 6, 'trace': /home/storage/Projects/Chips-Demo/demo/examples/radio/application.c : 18, 'op': 'return'}
  end

  
  always @(posedge clk)
  begin
    load_data <= memory[load_address];
    if(store_enable && state == execute) begin
      memory[store_address] <= store_data;
    end
  end


  //////////////////////////////////////////////////////////////////////////////
  // PIPELINE STAGE 1 -- FETCH INSTRUCTION
  //                                                                            
  
  always @(posedge clk)
  begin
    //implement memory for instructions
    if (state == instruction_fetch || state == operand_fetch || state == execute) begin
      instruction <= instructions[program_counter];
      program_counter_1 <= program_counter;
    end
  end

  assign opcode    = instruction[28:24];
  assign address_z = instruction[23:20];
  assign address_a = instruction[19:16];
  assign address_b = instruction[3:0];
  assign literal   = instruction[15:0];

  //////////////////////////////////////////////////////////////////////////////
  // PIPELINE STAGE 2 -- FETCH OPERANDS
  //                                                                            
  
  always @(posedge clk)
  begin
    if (write_enable) begin
      registers[address_z_3] <= result;
    end
    if (state == operand_fetch || state == execute) begin
      opcode_2 <= opcode;
      literal_2 <= literal;
      address_a_2 <= address_a;
      address_b_2 <= address_b;
      address_z_2 <= address_z;
      program_counter_2 <= program_counter_1;
    end
  end
  assign register_a = registers[address_a_2];
  assign register_b = registers[address_b_2];
  assign operand_a = (address_a_2 == address_z_3 && write_enable)?result:register_a;
  assign operand_b = (address_b_2 == address_z_3 && write_enable)?result:register_b;
  assign store_address = operand_a;
  assign load_address = operand_a;
  assign store_data = operand_b;
  assign store_enable = (opcode_2==2);

  //////////////////////////////////////////////////////////////////////////////
  // PIPELINE STAGE 3 -- EXECUTE
  //                                                                            
  
  always @(posedge clk)
  begin

  write_enable <= 0;
  timer_clock <= timer_clock + 1;
  case(state)

    //instruction_fetch
    instruction_fetch: begin
      program_counter <= program_counter + 1;
      state <= operand_fetch;
    end
    //operand_fetch
    operand_fetch: begin
      program_counter <= program_counter + 1;
      state <= execute;
    end
    //execute
    execute: begin
      program_counter <= program_counter + 1;
      address_z_3 <= address_z_2;
      case(opcode_2)

        //literal
        16'd0:
        begin
          result<=$signed(literal_2);
          write_enable <= 1;
        end

        //addl
        16'd1:
        begin
          result<=operand_a + literal_2;
          write_enable <= 1;
        end

        //store
        16'd2:
        begin
        end

        //call
        16'd3:
        begin
          result <= program_counter_2 + 1;
          write_enable <= 1;
          program_counter <= literal_2;
          state <= instruction_fetch;
        end

        //stop
        16'd4:
        begin
        state <= stop;
        end

        //literal_hi
        16'd5:
        begin
          result<= {literal_2, operand_a[15:0]};
          write_enable <= 1;
        end

        //load
        16'd6:
        begin
          state <= load;
        end

        //write
        16'd7:
        begin
          state <= write;
          write_output <= operand_a;
          write_value <= operand_b;
        end

        //a_hi
        16'd8:
        begin
          a_hi <= operand_a;
          result <= a_hi;
          write_enable <= 1;
        end

        //a_lo
        16'd9:
        begin
          a_lo <= operand_a;
          result <= a_lo;
          write_enable <= 1;
        end

        //long_to_double
        16'd10:
        begin
          long_to_double_in <= {a_hi, a_lo};
          state <= long_to_double_write_a;
        end

        //b_hi
        16'd11:
        begin
          b_hi <= operand_a;
          result <= b_hi;
          write_enable <= 1;
        end

        //b_lo
        16'd12:
        begin
          b_lo <= operand_a;
          result <= b_lo;
          write_enable <= 1;
        end

        //long_float_divide
        16'd13:
        begin
          double_divider_a <= {a_hi, a_lo};
          double_divider_b <= {b_hi, b_lo};
          state <= double_divider_write_a;
        end

        //double_to_long
        16'd14:
        begin
          double_to_long_in <= {a_hi, a_lo};
          state <= double_to_long_write_a;
        end

        //read
        16'd15:
        begin
          state <= read;
          read_input <= operand_a;
        end

        //shift_right
        16'd16:
        begin
          if(operand_b < 32) begin
            result <= $signed(operand_a) >>> operand_b;
            carry <= operand_a << (32-operand_b);
          end else begin
            result <= operand_a[31]?-1:0;
            carry <= operand_a;
          end
          write_enable <= 1;
        end

        //subtract
        16'd17:
        begin
          long_result = operand_a + (~operand_b) + 1;
          result <= long_result[31:0];
          carry[0] <= ~long_result[32];
          write_enable <= 1;
        end

        //add
        16'd18:
        begin
          long_result = operand_a + operand_b;
          result <= long_result[31:0];
          carry[0] <= long_result[32];
          write_enable <= 1;
        end

        //greater
        16'd19:
        begin
          result <= $signed(operand_a) > $signed(operand_b);
          write_enable <= 1;
        end

        //jmp_if_false
        16'd20:
        begin
          if (operand_a == 0) begin
            program_counter <= literal_2;
            state <= instruction_fetch;
          end
        end

        //goto
        16'd21:
        begin
          program_counter <= literal_2;
          state <= instruction_fetch;
        end

        //return
        16'd22:
        begin
          program_counter <= operand_a;
          state <= instruction_fetch;
        end

        //equal
        16'd23:
        begin
          result <= operand_a == operand_b;
          write_enable <= 1;
        end

        //multiply
        16'd24:
        begin
          product_a <= operand_a[15:0]  * operand_b[15:0];
          product_b <= operand_a[15:0]  * operand_b[31:16];
          product_c <= operand_a[31:16] * operand_b[15:0];
          product_d <= operand_a[31:16] * operand_b[31:16];
          state <= multiply;
        end

        //greater_equal
        16'd25:
        begin
          result <= $signed(operand_a) >= $signed(operand_b);
          write_enable <= 1;
        end

      endcase

    end

    multiply:
    begin
      long_result = product_a +
                    (product_b << 16) +
                    (product_c << 16) +
                    (product_d << 32);
      result <= long_result[31:0];
      carry <= long_result[63:32];
      write_enable <= 1;
      state <= execute;
    end

    read:
    begin
      case(read_input)
      0:
      begin
        s_input_eth_in_ack <= 1;
        if (s_input_eth_in_ack && input_eth_in_stb) begin
          result <= input_eth_in;
          write_enable <= 1;
          s_input_eth_in_ack <= 0;
          state <= execute;
        end
      end
      1:
      begin
        s_input_audio_in_ack <= 1;
        if (s_input_audio_in_ack && input_audio_in_stb) begin
          result <= input_audio_in;
          write_enable <= 1;
          s_input_audio_in_ack <= 0;
          state <= execute;
        end
      end
      2:
      begin
        s_input_rs232_rx_ack <= 1;
        if (s_input_rs232_rx_ack && input_rs232_rx_stb) begin
          result <= input_rs232_rx;
          write_enable <= 1;
          s_input_rs232_rx_ack <= 0;
          state <= execute;
        end
      end
      endcase
    end

    write:
    begin
      case(write_output)
      3:
      begin
        s_output_eth_out_stb <= 1;
        s_output_eth_out <= write_value;
        if (output_eth_out_ack && s_output_eth_out_stb) begin
          s_output_eth_out_stb <= 0;
          state <= execute;
        end
      end
      4:
      begin
        s_output_audio_out_stb <= 1;
        s_output_audio_out <= write_value;
        if (output_audio_out_ack && s_output_audio_out_stb) begin
          s_output_audio_out_stb <= 0;
          state <= execute;
        end
      end
      5:
      begin
        s_output_frequency_out_stb <= 1;
        s_output_frequency_out <= write_value;
        if (output_frequency_out_ack && s_output_frequency_out_stb) begin
          s_output_frequency_out_stb <= 0;
          state <= execute;
        end
      end
      6:
      begin
        s_output_samples_out_stb <= 1;
        s_output_samples_out <= write_value;
        if (output_samples_out_ack && s_output_samples_out_stb) begin
          s_output_samples_out_stb <= 0;
          state <= execute;
        end
      end
      7:
      begin
        s_output_rs232_tx_stb <= 1;
        s_output_rs232_tx <= write_value;
        if (output_rs232_tx_ack && s_output_rs232_tx_stb) begin
          s_output_rs232_tx_stb <= 0;
          state <= execute;
        end
      end
      endcase
    end

    load:
    begin
        result <= load_data;
        write_enable <= 1;
        state <= execute;
    end

    wait_state:
    begin
      if (timer) begin
        timer <= timer - 1;
      end else begin
        state <= execute;
      end
    end

    stop:
    begin
    end

    double_divider_write_a:
    begin
      double_divider_a_stb <= 1;
      if (double_divider_a_stb && double_divider_a_ack) begin
        double_divider_a_stb <= 0;
        state <= double_divider_write_b;
      end
    end

    double_divider_write_b:
    begin
      double_divider_b_stb <= 1;
      if (double_divider_b_stb && double_divider_b_ack) begin
        double_divider_b_stb <= 0;
        state <= double_divider_read_z;
      end
    end

    double_divider_read_z:
    begin
      double_divider_z_ack <= 1;
      if (double_divider_z_stb && double_divider_z_ack) begin
        a_lo <= double_divider_z[31:0];
        a_hi <= double_divider_z[63:32];
        double_divider_z_ack <= 0;
        state <= execute;
      end
    end

     double_to_long_write_a:
     begin
       double_to_long_in_stb <= 1;
       if (double_to_long_in_stb && double_to_long_in_ack) begin
         double_to_long_in_stb <= 0;
         state <= double_to_long_read_z;
       end
     end

     double_to_long_read_z:
     begin
       double_to_long_out_ack <= 1;
       if (double_to_long_out_stb && double_to_long_out_ack) begin
         double_to_long_out_ack <= 0;
         a_lo <= double_to_long_out[31:0];
         a_hi <= double_to_long_out[63:32];
         state <= execute;
       end
     end

     long_to_double_write_a:
     begin
       long_to_double_in_stb <= 1;
       if (long_to_double_in_stb && long_to_double_in_ack) begin
         long_to_double_in_stb <= 0;
         state <= long_to_double_read_z;
       end
     end

     long_to_double_read_z:
     begin
       long_to_double_out_ack <= 1;
       if (long_to_double_out_stb && long_to_double_out_ack) begin
         long_to_double_out_ack <= 0;
         a_lo <= long_to_double_out[31:0];
         a_hi <= long_to_double_out[63:32];
         state <= execute;
       end
     end

    endcase

    if (rst == 1'b1) begin
      timer <= 0;
      timer_clock <= 0;
      program_counter <= 0;
      address_z_3 <= 0;
      result <= 0;
      a = 0;
      b = 0;
      z = 0;
      state <= instruction_fetch;
      s_input_eth_in_ack <= 0;
      s_input_audio_in_ack <= 0;
      s_input_rs232_rx_ack <= 0;
      s_output_eth_out_stb <= 0;
      s_output_audio_out_stb <= 0;
      s_output_frequency_out_stb <= 0;
      s_output_samples_out_stb <= 0;
      s_output_rs232_tx_stb <= 0;
      double_divider_a_stb <= 0;
      double_divider_b_stb <= 0;
      double_divider_z_ack <= 0;
      double_to_long_in_stb <= 0;
      double_to_long_out_ack <= 0;
      long_to_double_in_stb <= 0;
      long_to_double_out_ack <= 0;
    end
  end
  assign input_eth_in_ack = s_input_eth_in_ack;
  assign input_audio_in_ack = s_input_audio_in_ack;
  assign input_rs232_rx_ack = s_input_rs232_rx_ack;
  assign output_eth_out_stb = s_output_eth_out_stb;
  assign output_eth_out = s_output_eth_out;
  assign output_audio_out_stb = s_output_audio_out_stb;
  assign output_audio_out = s_output_audio_out;
  assign output_frequency_out_stb = s_output_frequency_out_stb;
  assign output_frequency_out = s_output_frequency_out;
  assign output_samples_out_stb = s_output_samples_out_stb;
  assign output_samples_out = s_output_samples_out;
  assign output_rs232_tx_stb = s_output_rs232_tx_stb;
  assign output_rs232_tx = s_output_rs232_tx;

endmodule
